-- WRPC LM32 RAM initialization: --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.memory_loader_pkg.all;
use work.genram_pkg.all;

package wrc_bin_pkg is
  constant c_wrc_bin_init : t_ram_fast_load ( 0 to 32767 ) := (
        0 => x"98000000",     1 => x"d0000000",     2 => x"d0200000",
        3 => x"78010000",     4 => x"38210000",     5 => x"d0e10000",
        6 => x"f800003a",     7 => x"34000000",     8 => x"00000000",
        9 => x"00000000",    10 => x"00000000",    11 => x"00000000",
       12 => x"00000000",    13 => x"00000000",    14 => x"00000000",
       15 => x"00000000",    16 => x"00000000",    17 => x"00000000",
       18 => x"00000000",    19 => x"00000000",    20 => x"00000000",
       21 => x"00000000",    22 => x"00000000",    23 => x"00000000",
       24 => x"00000000",    25 => x"00000000",    26 => x"00000000",
       27 => x"00000000",    28 => x"00000000",    29 => x"00000000",
       30 => x"00000000",    31 => x"00000000",    32 => x"57525043",
       33 => x"2d2d2d2d",    34 => x"01234567",    35 => x"89abcdef",
       36 => x"00018f4c",    37 => x"00000000",    38 => x"00016178",
       39 => x"00000000",    40 => x"00000000",    41 => x"00000000",
       42 => x"00000000",    43 => x"00000000",    44 => x"00000000",
       45 => x"00000000",    46 => x"00000000",    47 => x"00000000",
       48 => x"5b9d0000",    49 => x"f800001e",    50 => x"34010002",
       51 => x"f800462b",    52 => x"e000002e",    53 => x"34000000",
       54 => x"34000000",    55 => x"34000000",    56 => x"00000000",
       57 => x"00000000",    58 => x"00000000",    59 => x"00000000",
       60 => x"00000000",    61 => x"00000000",    62 => x"00000000",
       63 => x"00000000",    64 => x"98000000",    65 => x"781c0001",
       66 => x"3b9cfffc",    67 => x"78010001",    68 => x"38217578",
       69 => x"34020000",    70 => x"78030001",    71 => x"386392c8",
       72 => x"c8611800",    73 => x"f8004bf8",    74 => x"34010000",
       75 => x"34020000",    76 => x"34030000",    77 => x"f800010e",
       78 => x"e0000000",    79 => x"379cffc4",    80 => x"5b810004",
       81 => x"5b820008",    82 => x"5b83000c",    83 => x"5b840010",
       84 => x"5b850014",    85 => x"5b860018",    86 => x"5b87001c",
       87 => x"5b880020",    88 => x"5b890024",    89 => x"5b8a0028",
       90 => x"5b9e0034",    91 => x"5b9f0038",    92 => x"2b81003c",
       93 => x"5b810030",    94 => x"bb800800",    95 => x"3421003c",
       96 => x"5b81002c",    97 => x"c3a00000",    98 => x"2b810004",
       99 => x"2b820008",   100 => x"2b83000c",   101 => x"2b840010",
      102 => x"2b850014",   103 => x"2b860018",   104 => x"2b87001c",
      105 => x"2b880020",   106 => x"2b890024",   107 => x"2b8a0028",
      108 => x"2b9d0030",   109 => x"2b9e0034",   110 => x"2b9f0038",
      111 => x"2b9c002c",   112 => x"34000000",   113 => x"c3c00000",
      114 => x"90001000",   115 => x"3401fffe",   116 => x"a0410800",
      117 => x"d0010000",   118 => x"90201000",   119 => x"3401fffe",
      120 => x"a0410800",   121 => x"d0210000",   122 => x"c3a00000",
      123 => x"90001000",   124 => x"3401fffe",   125 => x"a0410800",
      126 => x"d0010000",   127 => x"90201000",   128 => x"38420001",
      129 => x"d0220000",   130 => x"38210001",   131 => x"d0010000",
      132 => x"c3a00000",   133 => x"379cfff0",   134 => x"5b8b0008",
      135 => x"5b9d0004",   136 => x"f80037e8",   137 => x"f8004183",
      138 => x"f8004179",   139 => x"78010001",   140 => x"382136d4",
      141 => x"f8003162",   142 => x"34010001",   143 => x"f800370e",
      144 => x"f8003f2a",   145 => x"78010001",   146 => x"382191d0",
      147 => x"58200000",   148 => x"f8003e50",   149 => x"f800391d",
      150 => x"34010000",   151 => x"f80034ee",   152 => x"34010000",
      153 => x"34020050",   154 => x"f8003b71",   155 => x"3782000c",
      156 => x"34010000",   157 => x"f8003de1",   158 => x"3402ffff",
      159 => x"5c220010",   160 => x"78010001",   161 => x"382136f0",
      162 => x"f800314d",   163 => x"34010022",   164 => x"3381000c",
      165 => x"34010033",   166 => x"3381000d",   167 => x"34010044",
      168 => x"3381000e",   169 => x"34010055",   170 => x"3381000f",
      171 => x"34010066",   172 => x"33810010",   173 => x"34010077",
      174 => x"33810011",   175 => x"4384000e",   176 => x"4385000f",
      177 => x"43860010",   178 => x"43870011",   179 => x"4383000d",
      180 => x"4382000c",   181 => x"78010001",   182 => x"38213714",
      183 => x"f8003138",   184 => x"378b000c",   185 => x"b9600800",
      186 => x"f8003304",   187 => x"b9600800",   188 => x"f8003924",
      189 => x"34020001",   190 => x"34010001",   191 => x"f8003251",
      192 => x"f8003564",   193 => x"f8003a3b",   194 => x"f800029f",
      195 => x"78020001",   196 => x"38426170",   197 => x"34010002",
      198 => x"f80038bb",   199 => x"f8004655",   200 => x"f800276c",
      201 => x"f8002043",   202 => x"78030001",   203 => x"38635a28",
      204 => x"78010001",   205 => x"28620000",   206 => x"38217578",
      207 => x"58200000",   208 => x"78010001",   209 => x"3821f800",
      210 => x"58220000",   211 => x"34010003",   212 => x"f80002eb",
      213 => x"f800029e",   214 => x"78020001",   215 => x"34010000",
      216 => x"38427580",   217 => x"f8003a72",   218 => x"2b9d0004",
      219 => x"2b8b0008",   220 => x"379c0010",   221 => x"c3a00000",
      222 => x"379cfff8",   223 => x"5b8b0008",   224 => x"5b9d0004",
      225 => x"34010000",   226 => x"f8003260",   227 => x"b8205800",
      228 => x"78010001",   229 => x"38216174",   230 => x"28240000",
      231 => x"7d620000",   232 => x"64830000",   233 => x"a0431800",
      234 => x"4460000d",   235 => x"78010001",   236 => x"382192a8",
      237 => x"28210000",   238 => x"34020002",   239 => x"58220004",
      240 => x"f800371a",   241 => x"f8000282",   242 => x"78010001",
      243 => x"382192a0",   244 => x"34020001",   245 => x"58220000",
      246 => x"e0000014",   247 => x"65610000",   248 => x"7c840000",
      249 => x"a0240800",   250 => x"44230012",   251 => x"78010001",
      252 => x"382192a8",   253 => x"28210000",   254 => x"34020002",
      255 => x"58220008",   256 => x"78010001",   257 => x"382192a0",
      258 => x"58220000",   259 => x"f8000296",   260 => x"34010002",
      261 => x"34020000",   262 => x"34030001",   263 => x"f8004620",
      264 => x"34010000",   265 => x"f8003a72",   266 => x"34010001",
      267 => x"e0000008",   268 => x"fc411000",   269 => x"78010001",
      270 => x"c8021000",   271 => x"382192a0",   272 => x"20420003",
      273 => x"58220000",   274 => x"34010000",   275 => x"78020001",
      276 => x"38426174",   277 => x"584b0000",   278 => x"2b9d0004",
      279 => x"2b8b0008",   280 => x"379c0008",   281 => x"c3a00000",
      282 => x"379cfffc",   283 => x"5b9d0004",   284 => x"f8003693",
      285 => x"78020001",   286 => x"78030001",   287 => x"38637584",
      288 => x"38427588",   289 => x"28640000",   290 => x"28450000",
      291 => x"58610000",   292 => x"340303e8",   293 => x"c8a42000",
      294 => x"b4812000",   295 => x"58440000",   296 => x"34010000",
      297 => x"50640009",   298 => x"78010000",   299 => x"382100a0",
      300 => x"3484fc18",   301 => x"58440000",   302 => x"28220000",
      303 => x"34420001",   304 => x"58220000",   305 => x"34010001",
      306 => x"2b9d0004",   307 => x"379c0004",   308 => x"c3a00000",
      309 => x"379cfffc",   310 => x"5b9d0004",   311 => x"f8003678",
      312 => x"78020001",   313 => x"38427584",   314 => x"58410000",
      315 => x"2b9d0004",   316 => x"379c0004",   317 => x"c3a00000",
      318 => x"379cfff8",   319 => x"5b8b0008",   320 => x"5b9d0004",
      321 => x"78010001",   322 => x"38217578",   323 => x"28220000",
      324 => x"34010001",   325 => x"5c41000f",   326 => x"f8001d5f",
      327 => x"b8205800",   328 => x"f80040ea",   329 => x"3402001b",
      330 => x"44220005",   331 => x"78020001",   332 => x"38426168",
      333 => x"28410000",   334 => x"5c200008",   335 => x"f8001fbd",
      336 => x"78020001",   337 => x"38427578",   338 => x"58400000",
      339 => x"e0000003",   340 => x"f8001fc2",   341 => x"b8205800",
      342 => x"b9600800",   343 => x"2b9d0004",   344 => x"2b8b0008",
      345 => x"379c0008",   346 => x"c3a00000",   347 => x"379cffe0",
      348 => x"5b8b001c",   349 => x"5b8c0018",   350 => x"5b8d0014",
      351 => x"5b8e0010",   352 => x"5b8f000c",   353 => x"5b900008",
      354 => x"5b9d0004",   355 => x"780b0001",   356 => x"780c0001",
      357 => x"f800487d",   358 => x"396b7424",   359 => x"398c7574",
      360 => x"e0000005",   361 => x"29610008",   362 => x"44200002",
      363 => x"d8200000",   364 => x"356b001c",   365 => x"558bfffc",
      366 => x"780b0001",   367 => x"78010001",   368 => x"396b7424",
      369 => x"780f0001",   370 => x"780d0001",   371 => x"38215a2c",
      372 => x"39ef7574",   373 => x"39ad7580",   374 => x"282e0000",
      375 => x"b9608000",   376 => x"e0000025",   377 => x"2961000c",
      378 => x"5c200005",   379 => x"29610010",   380 => x"34210001",
      381 => x"59610010",   382 => x"e000000b",   383 => x"29620004",
      384 => x"44400003",   385 => x"28420000",   386 => x"44400007",
      387 => x"d8200000",   388 => x"29620010",   389 => x"b9606000",
      390 => x"b4411000",   391 => x"59620010",   392 => x"5c200002",
      393 => x"ba006000",   394 => x"34010000",   395 => x"37820020",
      396 => x"f80039bf",   397 => x"2b820020",   398 => x"29a10000",
      399 => x"c8410800",   400 => x"4c200002",   401 => x"b42e0800",
      402 => x"29830018",   403 => x"b4230800",   404 => x"59810018",
      405 => x"51c10006",   406 => x"c82e0800",   407 => x"59810018",
      408 => x"29810014",   409 => x"34210001",   410 => x"59810014",
      411 => x"59a20000",   412 => x"356b001c",   413 => x"55ebffdc",
      414 => x"f800482b",   415 => x"ba005800",   416 => x"e3fffffd",
      417 => x"379cffbc",   418 => x"5b8b0014",   419 => x"5b8c0010",
      420 => x"5b8d000c",   421 => x"5b8e0008",   422 => x"5b9d0004",
      423 => x"5b830030",   424 => x"78030001",   425 => x"3863758c",
      426 => x"5b82002c",   427 => x"5b840034",   428 => x"5b850038",
      429 => x"5b86003c",   430 => x"5b870040",   431 => x"5b880044",
      432 => x"286d0000",   433 => x"b8205800",   434 => x"b8407000",
      435 => x"34030000",   436 => x"44200002",   437 => x"28230018",
      438 => x"b86d1800",   439 => x"0063001c",   440 => x"4460001b",
      441 => x"780c0001",   442 => x"398c758c",   443 => x"39a10001",
      444 => x"59810000",   445 => x"29610028",   446 => x"37820018",
      447 => x"28230000",   448 => x"b9600800",   449 => x"d8600000",
      450 => x"78030001",   451 => x"38635a30",   452 => x"28620000",
      453 => x"2b81001c",   454 => x"598d0000",   455 => x"296b0334",
      456 => x"f800494d",   457 => x"780c0001",   458 => x"2b830018",
      459 => x"398c377c",   460 => x"b8202000",   461 => x"b9601000",
      462 => x"b9800800",   463 => x"f8003020",   464 => x"b9c00800",
      465 => x"37820030",   466 => x"f8002ffb",   467 => x"2b9d0004",
      468 => x"2b8b0014",   469 => x"2b8c0010",   470 => x"2b8d000c",
      471 => x"2b8e0008",   472 => x"379c0044",   473 => x"c3a00000",
      474 => x"379cfffc",   475 => x"5b9d0004",   476 => x"b8402800",
      477 => x"5c600005",   478 => x"78020001",   479 => x"38423798",
      480 => x"b8a01800",   481 => x"e000000c",   482 => x"34020001",
      483 => x"5c620006",   484 => x"78020001",   485 => x"384237b4",
      486 => x"b8a01800",   487 => x"28240008",   488 => x"e0000005",
      489 => x"28240004",   490 => x"78020001",   491 => x"384237cc",
      492 => x"b8a01800",   493 => x"fbffffb4",   494 => x"2b9d0004",
      495 => x"379c0004",   496 => x"c3a00000",   497 => x"379cffe8",
      498 => x"5b8b0018",   499 => x"5b8c0014",   500 => x"5b8d0010",
      501 => x"5b8e000c",   502 => x"5b9d0008",   503 => x"b8205800",
      504 => x"b8407000",   505 => x"b8606800",   506 => x"4460001a",
      507 => x"40480000",   508 => x"78020001",   509 => x"384267c4",
      510 => x"2108000f",   511 => x"3d030002",   512 => x"282600e4",
      513 => x"b4431000",   514 => x"28420000",   515 => x"282700e8",
      516 => x"78040001",   517 => x"5b820004",   518 => x"34030001",
      519 => x"34020005",   520 => x"388437e4",   521 => x"b9a02800",
      522 => x"f8000048",   523 => x"34010021",   524 => x"4c2d0006",
      525 => x"b9600800",   526 => x"b9c01000",   527 => x"b9a01800",
      528 => x"f8001607",   529 => x"44200003",   530 => x"340d0000",
      531 => x"340e0000",   532 => x"780c0001",   533 => x"29610000",
      534 => x"398c6654",   535 => x"e000002d",   536 => x"44410003",
      537 => x"358c000c",   538 => x"e000002a",   539 => x"59610004",
      540 => x"2961000c",   541 => x"59600008",   542 => x"44200006",
      543 => x"29820004",   544 => x"b9600800",   545 => x"34030000",
      546 => x"b9a02000",   547 => x"fbffffb7",   548 => x"29840008",
      549 => x"b9a01800",   550 => x"b9600800",   551 => x"b9c01000",
      552 => x"d8800000",   553 => x"b8201800",   554 => x"44200006",
      555 => x"29620334",   556 => x"29840004",   557 => x"78010001",
      558 => x"38213810",   559 => x"f8002fc0",   560 => x"29610004",
      561 => x"29630000",   562 => x"29820004",   563 => x"4461000a",
      564 => x"59610000",   565 => x"34010001",   566 => x"5961000c",
      567 => x"34030002",   568 => x"b9600800",   569 => x"34040000",
      570 => x"fbffffa0",   571 => x"34010000",   572 => x"e000000f",
      573 => x"b9600800",   574 => x"5960000c",   575 => x"34030001",
      576 => x"34040000",   577 => x"fbffff99",   578 => x"29610008",
      579 => x"e0000008",   580 => x"29820000",   581 => x"5c40ffd3",
      582 => x"29620334",   583 => x"78010001",   584 => x"3821382c",
      585 => x"f8002fa6",   586 => x"34012710",   587 => x"2b9d0008",
      588 => x"2b8b0018",   589 => x"2b8c0014",   590 => x"2b8d0010",
      591 => x"2b8e000c",   592 => x"379c0018",   593 => x"c3a00000",
      594 => x"379cffe4",   595 => x"5b8b0008",   596 => x"5b9d0004",
      597 => x"5b84000c",   598 => x"5b850010",   599 => x"b8805800",
      600 => x"5b860014",   601 => x"78040001",   602 => x"5b870018",
      603 => x"5b88001c",   604 => x"3884384c",   605 => x"34050000",
      606 => x"44200003",   607 => x"28240334",   608 => x"28250018",
      609 => x"78060001",   610 => x"38c6758c",   611 => x"28c10000",
      612 => x"3c420002",   613 => x"b8a12800",   614 => x"80a22800",
      615 => x"20a5000f",   616 => x"5465000c",   617 => x"78050001",
      618 => x"38a55af0",   619 => x"b4a22800",   620 => x"78060001",
      621 => x"28a20000",   622 => x"b8c00800",   623 => x"38213854",
      624 => x"f8002f7f",   625 => x"b9600800",   626 => x"37820010",
      627 => x"f8002f5a",   628 => x"2b9d0004",   629 => x"2b8b0008",
      630 => x"379c001c",   631 => x"c3a00000",   632 => x"379cfff8",
      633 => x"5b8b0008",   634 => x"5b9d0004",   635 => x"3402001c",
      636 => x"b8201800",   637 => x"340b0000",   638 => x"3405fffc",
      639 => x"34040003",   640 => x"e0000009",   641 => x"3421ffd0",
      642 => x"202600ff",   643 => x"50860002",   644 => x"e0000008",
      645 => x"bc220800",   646 => x"34630001",   647 => x"b9615800",
      648 => x"3442fffc",   649 => x"40610000",   650 => x"44200007",
      651 => x"5c45fff6",   652 => x"78010001",   653 => x"78020001",
      654 => x"38213860",   655 => x"38425ae0",   656 => x"f8002f5f",
      657 => x"b9600800",   658 => x"2b9d0004",   659 => x"2b8b0008",
      660 => x"379c0008",   661 => x"c3a00000",   662 => x"379cfffc",
      663 => x"5b9d0004",   664 => x"34030001",   665 => x"34010003",
      666 => x"34020000",   667 => x"f800448c",   668 => x"34010000",
      669 => x"34020001",   670 => x"f800461d",   671 => x"34010000",
      672 => x"2b9d0004",   673 => x"379c0004",   674 => x"c3a00000",
      675 => x"379cfff4",   676 => x"5b8b000c",   677 => x"5b8c0008",
      678 => x"5b9d0004",   679 => x"34010000",   680 => x"b8406000",
      681 => x"f8004548",   682 => x"45800005",   683 => x"642c0000",
      684 => x"c80c6000",   685 => x"398c0001",   686 => x"e000000f",
      687 => x"780b0001",   688 => x"396b7590",   689 => x"5c2c0004",
      690 => x"59600000",   691 => x"340cffff",   692 => x"e0000009",
      693 => x"29610000",   694 => x"340c0001",   695 => x"5c200006",
      696 => x"78020001",   697 => x"34010003",   698 => x"38426170",
      699 => x"f80036c6",   700 => x"596c0000",   701 => x"b9800800",
      702 => x"2b9d0004",   703 => x"2b8b000c",   704 => x"2b8c0008",
      705 => x"379c000c",   706 => x"c3a00000",   707 => x"34010000",
      708 => x"c3a00000",   709 => x"379cfffc",   710 => x"5b9d0004",
      711 => x"34010000",   712 => x"34020001",   713 => x"f80045f2",
      714 => x"34010000",   715 => x"2b9d0004",   716 => x"379c0004",
      717 => x"c3a00000",   718 => x"379cfffc",   719 => x"5b9d0004",
      720 => x"282102c8",   721 => x"28210010",   722 => x"2823000c",
      723 => x"44430004",   724 => x"5822000c",   725 => x"b8400800",
      726 => x"f80038a5",   727 => x"34010000",   728 => x"2b9d0004",
      729 => x"379c0004",   730 => x"c3a00000",   731 => x"379cfffc",
      732 => x"5b9d0004",   733 => x"f8003897",   734 => x"34020001",
      735 => x"5c200003",   736 => x"f80045cb",   737 => x"7c220000",
      738 => x"b8400800",   739 => x"2b9d0004",   740 => x"379c0004",
      741 => x"c3a00000",   742 => x"379cfff8",   743 => x"5b8b0008",
      744 => x"5b9d0004",   745 => x"b8202800",   746 => x"b8220800",
      747 => x"b8402000",   748 => x"b8605800",   749 => x"44200005",
      750 => x"34010001",   751 => x"b8a01000",   752 => x"b8801800",
      753 => x"f800381c",   754 => x"45600005",   755 => x"1562001f",
      756 => x"34010002",   757 => x"b9601800",   758 => x"f8003817",
      759 => x"34010000",   760 => x"2b9d0004",   761 => x"2b8b0008",
      762 => x"379c0008",   763 => x"c3a00000",   764 => x"379cfffc",
      765 => x"5b9d0004",   766 => x"b8201000",   767 => x"3401ffff",
      768 => x"f8004502",   769 => x"34010000",   770 => x"2b9d0004",
      771 => x"379c0004",   772 => x"c3a00000",   773 => x"379cff24",
      774 => x"5b8b0014",   775 => x"5b8c0010",   776 => x"5b8d000c",
      777 => x"5b8e0008",   778 => x"5b9d0004",   779 => x"b8406000",
      780 => x"28220330",   781 => x"b8807000",   782 => x"37810018",
      783 => x"b8605800",   784 => x"b8a06800",   785 => x"f8001d54",
      786 => x"45c00005",   787 => x"78010001",   788 => x"38216ffc",
      789 => x"28210000",   790 => x"59c10000",   791 => x"45a00003",
      792 => x"2b8100cc",   793 => x"59a10000",   794 => x"2b82006c",
      795 => x"3401fffd",   796 => x"44400013",   797 => x"45800007",
      798 => x"2b820060",   799 => x"2b810058",   800 => x"b4410800",
      801 => x"2b8200a0",   802 => x"b4220800",   803 => x"59810000",
      804 => x"2b820068",   805 => x"3401fffd",   806 => x"44400009",
      807 => x"34010000",   808 => x"45600007",   809 => x"2b830064",
      810 => x"2b82005c",   811 => x"b4621000",   812 => x"2b8300a4",
      813 => x"b4431000",   814 => x"59620000",   815 => x"2b9d0004",
      816 => x"2b8b0014",   817 => x"2b8c0010",   818 => x"2b8d000c",
      819 => x"2b8e0008",   820 => x"379c00dc",   821 => x"c3a00000",
      822 => x"34010000",   823 => x"c3a00000",   824 => x"34010000",
      825 => x"c3a00000",   826 => x"379cffec",   827 => x"5b8b000c",
      828 => x"5b8c0008",   829 => x"5b9d0004",   830 => x"34040000",
      831 => x"b8406000",   832 => x"b8605800",   833 => x"37820010",
      834 => x"37830014",   835 => x"34050000",   836 => x"5b800014",
      837 => x"5b800010",   838 => x"fbffffbf",   839 => x"34010001",
      840 => x"5d810003",   841 => x"2b810010",   842 => x"e0000002",
      843 => x"2b810014",   844 => x"59610000",   845 => x"34010001",
      846 => x"2b9d0004",   847 => x"2b8b000c",   848 => x"2b8c0008",
      849 => x"379c0014",   850 => x"c3a00000",   851 => x"379cfffc",
      852 => x"5b9d0004",   853 => x"f800302e",   854 => x"34010000",
      855 => x"2b9d0004",   856 => x"379c0004",   857 => x"c3a00000",
      858 => x"379cfffc",   859 => x"5b9d0004",   860 => x"f8003032",
      861 => x"34010000",   862 => x"2b9d0004",   863 => x"379c0004",
      864 => x"c3a00000",   865 => x"379cfffc",   866 => x"5b9d0004",
      867 => x"f800350d",   868 => x"f8003e9f",   869 => x"f8003ea7",
      870 => x"78010001",   871 => x"78020001",   872 => x"38423900",
      873 => x"382138d0",   874 => x"f8002e85",   875 => x"34010000",
      876 => x"2b9d0004",   877 => x"379c0004",   878 => x"c3a00000",
      879 => x"78010001",   880 => x"38217594",   881 => x"28210000",
      882 => x"c3a00000",   883 => x"379cfff8",   884 => x"5b8b0008",
      885 => x"5b9d0004",   886 => x"78010001",   887 => x"3821391c",
      888 => x"f8002e77",   889 => x"78010001",   890 => x"78020001",
      891 => x"38426824",   892 => x"382164ec",   893 => x"780b0001",
      894 => x"f800199c",   895 => x"396b6178",   896 => x"34030000",
      897 => x"b9600800",   898 => x"34020000",   899 => x"fbfffe6e",
      900 => x"78020001",   901 => x"38426530",   902 => x"58410000",
      903 => x"f8003428",   904 => x"78020001",   905 => x"3842759c",
      906 => x"58410000",   907 => x"296102c8",   908 => x"28210010",
      909 => x"58200068",   910 => x"b9600800",   911 => x"f8000ad5",
      912 => x"78010001",   913 => x"38217598",   914 => x"34020001",
      915 => x"58220000",   916 => x"34010000",   917 => x"2b9d0004",
      918 => x"2b8b0008",   919 => x"379c0008",   920 => x"c3a00000",
      921 => x"379cfff4",   922 => x"5b8b000c",   923 => x"5b8c0008",
      924 => x"5b9d0004",   925 => x"780b0001",   926 => x"396b6178",
      927 => x"296102c8",   928 => x"282c0010",   929 => x"78010001",
      930 => x"38213928",   931 => x"f8002e4c",   932 => x"29810000",
      933 => x"34020000",   934 => x"28230034",   935 => x"b9600800",
      936 => x"d8600000",   937 => x"78010001",   938 => x"34020000",
      939 => x"340301b8",   940 => x"59800040",   941 => x"31800035",
      942 => x"38216288",   943 => x"f8004892",   944 => x"78010001",
      945 => x"38217598",   946 => x"58200000",   947 => x"b9600800",
      948 => x"0d60010c",   949 => x"f8000aaf",   950 => x"78010001",
      951 => x"382164ec",   952 => x"f80019ab",   953 => x"34010000",
      954 => x"2b9d0004",   955 => x"2b8b000c",   956 => x"2b8c0008",
      957 => x"379c000c",   958 => x"c3a00000",   959 => x"379cffec",
      960 => x"5b8b0014",   961 => x"5b8c0010",   962 => x"5b8d000c",
      963 => x"5b8e0008",   964 => x"5b9d0004",   965 => x"780b0001",
      966 => x"396b6178",   967 => x"b8206000",   968 => x"296102c8",
      969 => x"282d0010",   970 => x"78010001",   971 => x"38217594",
      972 => x"58200000",   973 => x"fbffffcc",   974 => x"34010002",
      975 => x"45810016",   976 => x"34020003",   977 => x"45820026",
      978 => x"34010001",   979 => x"5d81002e",   980 => x"78010001",
      981 => x"31ac0004",   982 => x"38216824",   983 => x"340e0006",
      984 => x"316c001d",   985 => x"302e0000",   986 => x"34020000",
      987 => x"34010001",   988 => x"34030001",   989 => x"f800434a",
      990 => x"29610020",   991 => x"2821000c",   992 => x"302e000e",
      993 => x"b9600800",   994 => x"f80012ab",   995 => x"380bea60",
      996 => x"e000001e",   997 => x"34010001",   998 => x"31a10004",
      999 => x"3161001d",  1000 => x"78010001",  1001 => x"38216824",
     1002 => x"340effbb",  1003 => x"302e0000",  1004 => x"34020000",
     1005 => x"34010002",  1006 => x"34030001",  1007 => x"f8004338",
     1008 => x"29610020",  1009 => x"2821000c",  1010 => x"302e000e",
     1011 => x"b9600800",  1012 => x"f8001299",  1013 => x"340b0fa0",
     1014 => x"e000000c",  1015 => x"31a10004",  1016 => x"3161001d",
     1017 => x"78010001",  1018 => x"38216824",  1019 => x"3402ffff",
     1020 => x"30220000",  1021 => x"34030001",  1022 => x"34010003",
     1023 => x"34020000",  1024 => x"f8004327",  1025 => x"340b0000",
     1026 => x"f80033ad",  1027 => x"78020001",  1028 => x"b8207000",
     1029 => x"b8400800",  1030 => x"38213934",  1031 => x"f8002de8",
     1032 => x"29a20000",  1033 => x"780d0001",  1034 => x"39ad3950",
     1035 => x"28430034",  1036 => x"78020001",  1037 => x"b8400800",
     1038 => x"38216178",  1039 => x"34020000",  1040 => x"d8600000",
     1041 => x"e000000e",  1042 => x"f8004502",  1043 => x"340103e8",
     1044 => x"f80033a0",  1045 => x"f800339a",  1046 => x"c82e1000",
     1047 => x"51620006",  1048 => x"78010001",  1049 => x"38213940",
     1050 => x"f8002dd5",  1051 => x"340bff8c",  1052 => x"e0000008",
     1053 => x"b9a00800",  1054 => x"f8002dd1",  1055 => x"34010000",
     1056 => x"f80043d1",  1057 => x"5c200002",  1058 => x"5d61fff0",
     1059 => x"340b0000",  1060 => x"78010001",  1061 => x"38214d20",
     1062 => x"f8002dc9",  1063 => x"7d620000",  1064 => x"65810001",
     1065 => x"a0410800",  1066 => x"44200005",  1067 => x"78010001",
     1068 => x"38216824",  1069 => x"34020034",  1070 => x"30220000",
     1071 => x"78010001",  1072 => x"38217594",  1073 => x"582c0000",
     1074 => x"b9600800",  1075 => x"2b9d0004",  1076 => x"2b8b0014",
     1077 => x"2b8c0010",  1078 => x"2b8d000c",  1079 => x"2b8e0008",
     1080 => x"379c0014",  1081 => x"c3a00000",  1082 => x"379cffec",
     1083 => x"5b8b0014",  1084 => x"5b8c0010",  1085 => x"5b8d000c",
     1086 => x"5b8e0008",  1087 => x"5b9d0004",  1088 => x"78010001",
     1089 => x"38217598",  1090 => x"28210000",  1091 => x"340e0000",
     1092 => x"44200024",  1093 => x"780b0001",  1094 => x"396b6178",
     1095 => x"29610024",  1096 => x"29620038",  1097 => x"78040001",
     1098 => x"28250008",  1099 => x"3403007c",  1100 => x"b9600800",
     1101 => x"3884625c",  1102 => x"d8a00000",  1103 => x"b8201800",
     1104 => x"4c010005",  1105 => x"29610370",  1106 => x"34210001",
     1107 => x"59610370",  1108 => x"e000000c",  1109 => x"5c20000b",
     1110 => x"780d0001",  1111 => x"f8003358",  1112 => x"39ad759c",
     1113 => x"29a20000",  1114 => x"780c0001",  1115 => x"398c6530",
     1116 => x"c8220800",  1117 => x"29820000",  1118 => x"5441000a",
     1119 => x"e0000011",  1120 => x"78010001",  1121 => x"38216178",
     1122 => x"28220040",  1123 => x"fbfffd8e",  1124 => x"78020001",
     1125 => x"38426530",  1126 => x"58410000",  1127 => x"340e0001",
     1128 => x"b9c00800",  1129 => x"2b9d0004",  1130 => x"2b8b0014",
     1131 => x"2b8c0010",  1132 => x"2b8d000c",  1133 => x"2b8e0008",
     1134 => x"379c0014",  1135 => x"c3a00000",  1136 => x"f800333f",
     1137 => x"59a10000",  1138 => x"34020000",  1139 => x"b9600800",
     1140 => x"34030000",  1141 => x"fbfffd7c",  1142 => x"59810000",
     1143 => x"e3fffff0",  1144 => x"379cffe8",  1145 => x"5b9d0018",
     1146 => x"b8205000",  1147 => x"40610005",  1148 => x"40640000",
     1149 => x"40650001",  1150 => x"40660002",  1151 => x"40670003",
     1152 => x"40680004",  1153 => x"5b810004",  1154 => x"40610006",
     1155 => x"b8404800",  1156 => x"b9401000",  1157 => x"5b810008",
     1158 => x"40610007",  1159 => x"5b81000c",  1160 => x"40610008",
     1161 => x"5b810010",  1162 => x"40610009",  1163 => x"b9201800",
     1164 => x"5b810014",  1165 => x"78010001",  1166 => x"38213958",
     1167 => x"f8002d60",  1168 => x"2b9d0018",  1169 => x"379c0018",
     1170 => x"c3a00000",  1171 => x"379cffd0",  1172 => x"5b8b0030",
     1173 => x"5b8c002c",  1174 => x"5b8d0028",  1175 => x"5b8e0024",
     1176 => x"5b8f0020",  1177 => x"5b90001c",  1178 => x"5b910018",
     1179 => x"5b920014",  1180 => x"5b930010",  1181 => x"5b94000c",
     1182 => x"5b950008",  1183 => x"5b9d0004",  1184 => x"b8603000",
     1185 => x"b8209800",  1186 => x"b8409000",  1187 => x"78010001",
     1188 => x"b880a800",  1189 => x"38213990",  1190 => x"ba601000",
     1191 => x"ba401800",  1192 => x"b8c02000",  1193 => x"b8a0a000",
     1194 => x"78110001",  1195 => x"f8002d44",  1196 => x"78100001",
     1197 => x"780f0001",  1198 => x"780e0001",  1199 => x"780d0001",
     1200 => x"b8205800",  1201 => x"340c0000",  1202 => x"3a3139a4",
     1203 => x"3a1039ac",  1204 => x"39ef4e44",  1205 => x"39ce4d20",
     1206 => x"39ad4ba0",  1207 => x"e0000017",  1208 => x"5cc00006",
     1209 => x"ba200800",  1210 => x"ba601000",  1211 => x"ba401800",
     1212 => x"f8002d33",  1213 => x"b5615800",  1214 => x"b6ac1000",
     1215 => x"40420000",  1216 => x"ba000800",  1217 => x"358c0001",
     1218 => x"f8002d2d",  1219 => x"21820003",  1220 => x"b42b5800",
     1221 => x"b9e03000",  1222 => x"5c400005",  1223 => x"2181000f",
     1224 => x"b9c03000",  1225 => x"44220002",  1226 => x"b9a03000",
     1227 => x"b8c00800",  1228 => x"f8002d23",  1229 => x"b5615800",
     1230 => x"2186000f",  1231 => x"4a8cffe9",  1232 => x"44c00005",
     1233 => x"78010001",  1234 => x"38214d20",  1235 => x"f8002d1c",
     1236 => x"b42b5800",  1237 => x"b9600800",  1238 => x"2b9d0004",
     1239 => x"2b8b0030",  1240 => x"2b8c002c",  1241 => x"2b8d0028",
     1242 => x"2b8e0024",  1243 => x"2b8f0020",  1244 => x"2b90001c",
     1245 => x"2b910018",  1246 => x"2b920014",  1247 => x"2b930010",
     1248 => x"2b94000c",  1249 => x"2b950008",  1250 => x"379c0030",
     1251 => x"c3a00000",  1252 => x"379cffb8",  1253 => x"5b8b0048",
     1254 => x"5b8c0044",  1255 => x"5b8d0040",  1256 => x"5b8e003c",
     1257 => x"5b8f0038",  1258 => x"5b900034",  1259 => x"5b910030",
     1260 => x"5b92002c",  1261 => x"5b930028",  1262 => x"5b940024",
     1263 => x"5b950020",  1264 => x"5b96001c",  1265 => x"5b970018",
     1266 => x"5b980014",  1267 => x"5b9d0010",  1268 => x"b8608000",
     1269 => x"40430001",  1270 => x"b8206000",  1271 => x"34010002",
     1272 => x"2063000f",  1273 => x"b8406800",  1274 => x"404e0000",
     1275 => x"44610006",  1276 => x"78010001",  1277 => x"b9801000",
     1278 => x"382139b4",  1279 => x"f8002cf0",  1280 => x"e000013f",
     1281 => x"40450002",  1282 => x"40460003",  1283 => x"21ce000f",
     1284 => x"3ca50008",  1285 => x"78010001",  1286 => x"b8c52800",
     1287 => x"41a60004",  1288 => x"34030002",  1289 => x"b9c02000",
     1290 => x"344b0022",  1291 => x"382139d4",  1292 => x"b9801000",
     1293 => x"f8002ce2",  1294 => x"41a2000c",  1295 => x"41a1000d",
     1296 => x"41a4000e",  1297 => x"41a30006",  1298 => x"3c420018",
     1299 => x"3c210010",  1300 => x"41a60007",  1301 => x"41a5000f",
     1302 => x"3c840008",  1303 => x"b8220800",  1304 => x"3c630008",
     1305 => x"b8812000",  1306 => x"78010001",  1307 => x"b8c31800",
     1308 => x"b8a42000",  1309 => x"b9801000",  1310 => x"38213a00",
     1311 => x"f8002cd0",  1312 => x"78020001",  1313 => x"b9800800",
     1314 => x"38423a24",  1315 => x"35a30014",  1316 => x"fbffff54",
     1317 => x"41a3001e",  1318 => x"41a4001f",  1319 => x"41a50021",
     1320 => x"3c630008",  1321 => x"78010001",  1322 => x"b8831800",
     1323 => x"41a40020",  1324 => x"38213a2c",  1325 => x"b9801000",
     1326 => x"f8002cc1",  1327 => x"3401000c",  1328 => x"55c100d1",
     1329 => x"78010001",  1330 => x"3dce0002",  1331 => x"38215b10",
     1332 => x"b42e0800",  1333 => x"28210000",  1334 => x"c0200000",
     1335 => x"78010001",  1336 => x"b9801000",  1337 => x"38213a58",
     1338 => x"f8002cb5",  1339 => x"41620002",  1340 => x"41610003",
     1341 => x"41640004",  1342 => x"3c420018",  1343 => x"3c210010",
     1344 => x"3c840008",  1345 => x"b8220800",  1346 => x"b8812000",
     1347 => x"41620006",  1348 => x"41610007",  1349 => x"41650008",
     1350 => x"3c420018",  1351 => x"3c210010",  1352 => x"3ca50008",
     1353 => x"b8220800",  1354 => x"b8a12800",  1355 => x"78030001",
     1356 => x"78010001",  1357 => x"41670005",  1358 => x"41660009",
     1359 => x"38213a70",  1360 => x"b9801000",  1361 => x"38633a80",
     1362 => x"e000001c",  1363 => x"78010001",  1364 => x"b9801000",
     1365 => x"38213a8c",  1366 => x"f8002c99",  1367 => x"41620002",
     1368 => x"41610003",  1369 => x"41640004",  1370 => x"3c420018",
     1371 => x"3c210010",  1372 => x"3c840008",  1373 => x"b8220800",
     1374 => x"b8812000",  1375 => x"41620006",  1376 => x"41610007",
     1377 => x"41650008",  1378 => x"3c420018",  1379 => x"3c210010",
     1380 => x"3ca50008",  1381 => x"b8220800",  1382 => x"41670005",
     1383 => x"41660009",  1384 => x"b8a12800",  1385 => x"78030001",
     1386 => x"78010001",  1387 => x"38213a70",  1388 => x"b9801000",
     1389 => x"38633aa8",  1390 => x"b8e42000",  1391 => x"b8c52800",
     1392 => x"f8002c7f",  1393 => x"e000008e",  1394 => x"78010001",
     1395 => x"b9801000",  1396 => x"38213ab8",  1397 => x"f8002c7a",
     1398 => x"41620002",  1399 => x"41610003",  1400 => x"41640004",
     1401 => x"3c420018",  1402 => x"3c210010",  1403 => x"3c840008",
     1404 => x"b8220800",  1405 => x"b8812000",  1406 => x"41620006",
     1407 => x"41610007",  1408 => x"41650008",  1409 => x"3c420018",
     1410 => x"3c210010",  1411 => x"3ca50008",  1412 => x"b8220800",
     1413 => x"b8a12800",  1414 => x"78030001",  1415 => x"78010001",
     1416 => x"41670005",  1417 => x"41660009",  1418 => x"38213a70",
     1419 => x"b9801000",  1420 => x"38633ad4",  1421 => x"e3ffffe1",
     1422 => x"78010001",  1423 => x"b9801000",  1424 => x"38213ae4",
     1425 => x"f8002c5e",  1426 => x"41620002",  1427 => x"41610003",
     1428 => x"41640004",  1429 => x"3c420018",  1430 => x"3c210010",
     1431 => x"3c840008",  1432 => x"b8220800",  1433 => x"b8812000",
     1434 => x"41620006",  1435 => x"41610007",  1436 => x"41650008",
     1437 => x"3c420018",  1438 => x"3c210010",  1439 => x"41670005",
     1440 => x"41660009",  1441 => x"3ca50008",  1442 => x"b8220800",
     1443 => x"780e0001",  1444 => x"39ce3b00",  1445 => x"b8a12800",
     1446 => x"78010001",  1447 => x"b9801000",  1448 => x"b9c01800",
     1449 => x"b8e42000",  1450 => x"b8c52800",  1451 => x"38213a70",
     1452 => x"f8002c43",  1453 => x"3563000a",  1454 => x"b9800800",
     1455 => x"b9c01000",  1456 => x"fbfffec8",  1457 => x"340b0036",
     1458 => x"e0000080",  1459 => x"78010001",  1460 => x"b9801000",
     1461 => x"38213b14",  1462 => x"f8002c39",  1463 => x"41620002",
     1464 => x"41610003",  1465 => x"41640004",  1466 => x"3c420018",
     1467 => x"3c210010",  1468 => x"3c840008",  1469 => x"b8220800",
     1470 => x"b8812000",  1471 => x"41620006",  1472 => x"41610007",
     1473 => x"41650008",  1474 => x"3c420018",  1475 => x"3c210010",
     1476 => x"41670005",  1477 => x"41660009",  1478 => x"3ca50008",
     1479 => x"b8220800",  1480 => x"b8a12800",  1481 => x"78030001",
     1482 => x"78010001",  1483 => x"b8e42000",  1484 => x"b8c52800",
     1485 => x"b9801000",  1486 => x"38633b30",  1487 => x"38213a70",
     1488 => x"f8002c1f",  1489 => x"41660010",  1490 => x"41670011",
     1491 => x"4165000f",  1492 => x"4164000e",  1493 => x"3cc60008",
     1494 => x"78010001",  1495 => x"78030001",  1496 => x"b8e63000",
     1497 => x"b9801000",  1498 => x"38633b5c",  1499 => x"38213b48",
     1500 => x"f8002c13",  1501 => x"4163000d",  1502 => x"41640012",
     1503 => x"78010001",  1504 => x"b9801000",  1505 => x"38213b80",
     1506 => x"f8002c0d",  1507 => x"41610018",  1508 => x"41640013",
     1509 => x"41650014",  1510 => x"41660015",  1511 => x"41670016",
     1512 => x"41680017",  1513 => x"5b810004",  1514 => x"41610019",
     1515 => x"78030001",  1516 => x"b9801000",  1517 => x"5b810008",
     1518 => x"4161001a",  1519 => x"38633bd8",  1520 => x"340b0040",
     1521 => x"5b81000c",  1522 => x"78010001",  1523 => x"38213ba8",
     1524 => x"f8002bfb",  1525 => x"e000003d",  1526 => x"78010001",
     1527 => x"b9801000",  1528 => x"38213bf8",  1529 => x"f8002bf6",
     1530 => x"78020001",  1531 => x"b9800800",  1532 => x"38423c14",
     1533 => x"b9601800",  1534 => x"fbfffe7a",  1535 => x"340b002c",
     1536 => x"e0000032",  1537 => x"340b0022",  1538 => x"e0000030",
     1539 => x"55f70009",  1540 => x"78010001",  1541 => x"b9801000",
     1542 => x"ba001800",  1543 => x"b9602000",  1544 => x"b9e02800",
     1545 => x"38213c30",  1546 => x"f8002be5",  1547 => x"e0000034",
     1548 => x"b5ab7000",  1549 => x"41d60002",  1550 => x"41c10003",
     1551 => x"41c30000",  1552 => x"3ed60008",  1553 => x"41c40001",
     1554 => x"b836b000",  1555 => x"41c10008",  1556 => x"41c50004",
     1557 => x"41c60005",  1558 => x"41c70006",  1559 => x"41c80007",
     1560 => x"5b810004",  1561 => x"41c10009",  1562 => x"3c630008",
     1563 => x"36d10004",  1564 => x"5b810008",  1565 => x"b8831800",
     1566 => x"baa00800",  1567 => x"b9801000",  1568 => x"ba202000",
     1569 => x"f8002bce",  1570 => x"4df10007",  1571 => x"ba400800",
     1572 => x"b9801000",  1573 => x"ba201800",  1574 => x"b9e02000",
     1575 => x"f8002bc8",  1576 => x"e0000008",  1577 => x"b9800800",
     1578 => x"ba801000",  1579 => x"ba601800",  1580 => x"35c4000a",
     1581 => x"36c5fffa",  1582 => x"fbfffe65",  1583 => x"ba207800",
     1584 => x"b56f5800",  1585 => x"e000000b",  1586 => x"78150001",
     1587 => x"78140001",  1588 => x"78130001",  1589 => x"78120001",
     1590 => x"34180002",  1591 => x"34170009",  1592 => x"3ab53c54",
     1593 => x"3a943cc0",  1594 => x"3a733cc8",  1595 => x"3a523c94",
     1596 => x"4d700003",  1597 => x"ca0b7800",  1598 => x"49f8ffc5",
     1599 => x"78020001",  1600 => x"78030001",  1601 => x"b9800800",
     1602 => x"38423cd4",  1603 => x"38633cdc",  1604 => x"b9a02000",
     1605 => x"ba002800",  1606 => x"fbfffe4d",  1607 => x"2b9d0010",
     1608 => x"2b8b0048",  1609 => x"2b8c0044",  1610 => x"2b8d0040",
     1611 => x"2b8e003c",  1612 => x"2b8f0038",  1613 => x"2b900034",
     1614 => x"2b910030",  1615 => x"2b92002c",  1616 => x"2b930028",
     1617 => x"2b940024",  1618 => x"2b950020",  1619 => x"2b96001c",
     1620 => x"2b970018",  1621 => x"2b980014",  1622 => x"379c0048",
     1623 => x"c3a00000",  1624 => x"379cfff0",  1625 => x"5b8b0010",
     1626 => x"5b8c000c",  1627 => x"5b8d0008",  1628 => x"5b9d0004",
     1629 => x"b8205800",  1630 => x"b8406800",  1631 => x"b8606000",
     1632 => x"4480000f",  1633 => x"2881000c",  1634 => x"78070001",
     1635 => x"28850000",  1636 => x"28860004",  1637 => x"38e75a24",
     1638 => x"5c200003",  1639 => x"78070001",  1640 => x"38e73ce4",
     1641 => x"78010001",  1642 => x"38213cf0",  1643 => x"b9601000",
     1644 => x"b8a01800",  1645 => x"b8a02000",  1646 => x"f8002b81",
     1647 => x"b9600800",  1648 => x"b9a01000",  1649 => x"b9801800",
     1650 => x"fbfffe72",  1651 => x"34010000",  1652 => x"2b9d0004",
     1653 => x"2b8b0010",  1654 => x"2b8c000c",  1655 => x"2b8d0008",
     1656 => x"379c0010",  1657 => x"c3a00000",  1658 => x"379cffe8",
     1659 => x"5b8b0018",  1660 => x"5b8c0014",  1661 => x"5b8d0010",
     1662 => x"5b8e000c",  1663 => x"5b8f0008",  1664 => x"5b9d0004",
     1665 => x"282d0000",  1666 => x"b8207800",  1667 => x"282e0004",
     1668 => x"b8406000",  1669 => x"340b0000",  1670 => x"34010000",
     1671 => x"34040000",  1672 => x"544d0006",  1673 => x"b9a00800",
     1674 => x"f80044d8",  1675 => x"882c1000",  1676 => x"b9602000",
     1677 => x"c9a26800",  1678 => x"34030000",  1679 => x"34020001",
     1680 => x"e000000b",  1681 => x"3d850001",  1682 => x"3d6b0001",
     1683 => x"f5856000",  1684 => x"3c630001",  1685 => x"b58b5800",
     1686 => x"b8a06000",  1687 => x"3c450001",  1688 => x"f4451000",
     1689 => x"b4431800",  1690 => x"b8a01000",  1691 => x"1565001f",
     1692 => x"c8ac3000",  1693 => x"f4c53000",  1694 => x"c8ab2800",
     1695 => x"c8a62800",  1696 => x"00a5001f",  1697 => x"34060001",
     1698 => x"55ab0004",  1699 => x"5dab0002",  1700 => x"55cc0002",
     1701 => x"34060000",  1702 => x"a0a63000",  1703 => x"5cc0ffea",
     1704 => x"556d000d",  1705 => x"5d6d0002",  1706 => x"558e000b",
     1707 => x"c9cc2800",  1708 => x"f4ae7000",  1709 => x"c9ab6800",
     1710 => x"c9ae6800",  1711 => x"b8a07000",  1712 => x"b4822800",
     1713 => x"f4852000",  1714 => x"b4230800",  1715 => x"b4810800",
     1716 => x"b8a02000",  1717 => x"3c65001f",  1718 => x"00420001",
     1719 => x"00630001",  1720 => x"b8a21000",  1721 => x"b8622800",
     1722 => x"44a00006",  1723 => x"3d65001f",  1724 => x"018c0001",
     1725 => x"016b0001",  1726 => x"b8ac6000",  1727 => x"e3ffffe9",
     1728 => x"59e10000",  1729 => x"b9c00800",  1730 => x"59e40004",
     1731 => x"2b9d0004",  1732 => x"2b8b0018",  1733 => x"2b8c0014",
     1734 => x"2b8d0010",  1735 => x"2b8e000c",  1736 => x"2b8f0008",
     1737 => x"379c0018",  1738 => x"c3a00000",  1739 => x"379cfff8",
     1740 => x"5b8b0008",  1741 => x"5b9d0004",  1742 => x"b8405800",
     1743 => x"f80030e0",  1744 => x"b42b0800",  1745 => x"5c200002",
     1746 => x"34010001",  1747 => x"2b9d0004",  1748 => x"2b8b0008",
     1749 => x"379c0008",  1750 => x"c3a00000",  1751 => x"379cfff8",
     1752 => x"5b8b0008",  1753 => x"5b9d0004",  1754 => x"78040001",
     1755 => x"b8405800",  1756 => x"78050001",  1757 => x"34020006",
     1758 => x"34030001",  1759 => x"38843dbc",  1760 => x"38a55b44",
     1761 => x"b9603000",  1762 => x"fbfffb70",  1763 => x"45600005",
     1764 => x"1562001f",  1765 => x"34010002",  1766 => x"b9601800",
     1767 => x"f8003426",  1768 => x"34010000",  1769 => x"2b9d0004",
     1770 => x"2b8b0008",  1771 => x"379c0008",  1772 => x"c3a00000",
     1773 => x"379cfff4",  1774 => x"5b8b000c",  1775 => x"5b8c0008",
     1776 => x"5b9d0004",  1777 => x"b8206000",  1778 => x"b8405800",
     1779 => x"b8603000",  1780 => x"44600008",  1781 => x"78040001",
     1782 => x"78050001",  1783 => x"34020006",  1784 => x"34030001",
     1785 => x"38843dc8",  1786 => x"38a55b64",  1787 => x"fbfffb57",
     1788 => x"b9800800",  1789 => x"b9601000",  1790 => x"fbffffd9",
     1791 => x"2b9d0004",  1792 => x"2b8b000c",  1793 => x"2b8c0008",
     1794 => x"379c000c",  1795 => x"c3a00000",  1796 => x"379cfff0",
     1797 => x"5b8b0010",  1798 => x"5b8c000c",  1799 => x"5b8d0008",
     1800 => x"5b9d0004",  1801 => x"b8206800",  1802 => x"44400012",
     1803 => x"284b0000",  1804 => x"284c0004",  1805 => x"34040003",
     1806 => x"1561001f",  1807 => x"b9601000",  1808 => x"b9801800",
     1809 => x"f800341a",  1810 => x"78040001",  1811 => x"78050001",
     1812 => x"b9a00800",  1813 => x"34020006",  1814 => x"34030001",
     1815 => x"38843df4",  1816 => x"38a55b78",  1817 => x"b9603000",
     1818 => x"b9803800",  1819 => x"fbfffb37",  1820 => x"34010000",
     1821 => x"2b9d0004",  1822 => x"2b8b0010",  1823 => x"2b8c000c",
     1824 => x"2b8d0008",  1825 => x"379c0010",  1826 => x"c3a00000",
     1827 => x"379cffe8",  1828 => x"5b8b000c",  1829 => x"5b8c0008",
     1830 => x"5b9d0004",  1831 => x"b8405800",  1832 => x"b8206000",
     1833 => x"37820018",  1834 => x"37810010",  1835 => x"f8003420",
     1836 => x"78020001",  1837 => x"3842758c",  1838 => x"2b860014",
     1839 => x"2b870018",  1840 => x"28410000",  1841 => x"59660000",
     1842 => x"59670004",  1843 => x"20210001",  1844 => x"5c200009",
     1845 => x"78040001",  1846 => x"78050001",  1847 => x"b9800800",
     1848 => x"34020006",  1849 => x"34030002",  1850 => x"38843df4",
     1851 => x"38a55b88",  1852 => x"fbfffb16",  1853 => x"34010000",
     1854 => x"2b9d0004",  1855 => x"2b8b000c",  1856 => x"2b8c0008",
     1857 => x"379c0018",  1858 => x"c3a00000",  1859 => x"379cffb0",
     1860 => x"5b8b001c",  1861 => x"5b8c0018",  1862 => x"5b8d0014",
     1863 => x"5b8e0010",  1864 => x"5b8f000c",  1865 => x"5b900008",
     1866 => x"5b9d0004",  1867 => x"28300058",  1868 => x"378c0040",
     1869 => x"b8407800",  1870 => x"b8206800",  1871 => x"78020001",
     1872 => x"340188f7",  1873 => x"b8607000",  1874 => x"0f81004c",
     1875 => x"38425ad8",  1876 => x"b9800800",  1877 => x"34030006",
     1878 => x"b8805800",  1879 => x"f800446c",  1880 => x"b9801000",
     1881 => x"ba000800",  1882 => x"b9e01800",  1883 => x"b9c02000",
     1884 => x"37850020",  1885 => x"f80022ef",  1886 => x"b8206000",
     1887 => x"45600011",  1888 => x"2b81003c",  1889 => x"2b870024",
     1890 => x"2b880028",  1891 => x"78040001",  1892 => x"78050001",
     1893 => x"5961000c",  1894 => x"59670000",  1895 => x"59680004",
     1896 => x"59600008",  1897 => x"b9a00800",  1898 => x"34020005",
     1899 => x"34030002",  1900 => x"38843e04",  1901 => x"38a55b98",
     1902 => x"b9803000",  1903 => x"fbfffae3",  1904 => x"4c0c0010",
     1905 => x"78010001",  1906 => x"3821758c",  1907 => x"28220000",
     1908 => x"29a10018",  1909 => x"b8410800",  1910 => x"00210014",
     1911 => x"34020001",  1912 => x"2021000f",  1913 => x"50410007",
     1914 => x"78010001",  1915 => x"38213e24",  1916 => x"b9e01000",
     1917 => x"b9c01800",  1918 => x"b9602000",  1919 => x"fbfffed9",
     1920 => x"b9800800",  1921 => x"2b9d0004",  1922 => x"2b8b001c",
     1923 => x"2b8c0018",  1924 => x"2b8d0014",  1925 => x"2b8e0010",
     1926 => x"2b8f000c",  1927 => x"2b900008",  1928 => x"379c0050",
     1929 => x"c3a00000",  1930 => x"379cffb8",  1931 => x"5b8b0014",
     1932 => x"5b8c0010",  1933 => x"5b8d000c",  1934 => x"5b8e0008",
     1935 => x"5b9d0004",  1936 => x"b8207000",  1937 => x"28210058",
     1938 => x"b8602800",  1939 => x"b8406800",  1940 => x"b8805800",
     1941 => x"37820038",  1942 => x"b8a02000",  1943 => x"b9a01800",
     1944 => x"37850018",  1945 => x"f8002241",  1946 => x"b8206000",
     1947 => x"4560000b",  1948 => x"2b81001c",  1949 => x"59610000",
     1950 => x"2b810020",  1951 => x"59610004",  1952 => x"2b810024",
     1953 => x"59610008",  1954 => x"2b810034",  1955 => x"5961000c",
     1956 => x"2b810030",  1957 => x"59610010",  1958 => x"4c0c0010",
     1959 => x"78040001",  1960 => x"3884758c",  1961 => x"28820000",
     1962 => x"29c10018",  1963 => x"b8410800",  1964 => x"00210014",
     1965 => x"34020001",  1966 => x"2021000f",  1967 => x"50410007",
     1968 => x"78010001",  1969 => x"38213e2c",  1970 => x"b9a01000",
     1971 => x"b9801800",  1972 => x"b9602000",  1973 => x"fbfffea3",
     1974 => x"b9800800",  1975 => x"2b9d0004",  1976 => x"2b8b0014",
     1977 => x"2b8c0010",  1978 => x"2b8d000c",  1979 => x"2b8e0008",
     1980 => x"379c0048",  1981 => x"c3a00000",  1982 => x"379cfffc",
     1983 => x"5b9d0004",  1984 => x"28210058",  1985 => x"f80021bf",
     1986 => x"34010000",  1987 => x"2b9d0004",  1988 => x"379c0004",
     1989 => x"c3a00000",  1990 => x"379cffd4",  1991 => x"5b8b0010",
     1992 => x"5b8c000c",  1993 => x"5b8d0008",  1994 => x"5b9d0004",
     1995 => x"b8205800",  1996 => x"28210058",  1997 => x"44200002",
     1998 => x"f80021b2",  1999 => x"b9600800",  2000 => x"f8000d2a",
     2001 => x"378c0014",  2002 => x"340188f7",  2003 => x"78020001",
     2004 => x"0f810020",  2005 => x"38425ad8",  2006 => x"b9800800",
     2007 => x"34030006",  2008 => x"f80043eb",  2009 => x"78010001",
     2010 => x"b9801000",  2011 => x"38216620",  2012 => x"34030001",
     2013 => x"34040000",  2014 => x"f8002159",  2015 => x"b8206000",
     2016 => x"4420000e",  2017 => x"378d0028",  2018 => x"b9a01000",
     2019 => x"f8002143",  2020 => x"b9a01000",  2021 => x"34030006",
     2022 => x"35610060",  2023 => x"f80043dc",  2024 => x"3561004c",
     2025 => x"596c0058",  2026 => x"b9a01000",  2027 => x"34030006",
     2028 => x"f80043d7",  2029 => x"596c0044",  2030 => x"34010000",
     2031 => x"2b9d0004",  2032 => x"2b8b0010",  2033 => x"2b8c000c",
     2034 => x"2b8d0008",  2035 => x"379c002c",  2036 => x"c3a00000",
     2037 => x"379cfff8",  2038 => x"5b8b0008",  2039 => x"5b9d0004",
     2040 => x"78040001",  2041 => x"78050001",  2042 => x"34020002",
     2043 => x"34030002",  2044 => x"38843f18",  2045 => x"38a55bf8",
     2046 => x"b8205800",  2047 => x"fbfffa53",  2048 => x"296302c8",
     2049 => x"28610010",  2050 => x"28220064",  2051 => x"34010000",
     2052 => x"44400010",  2053 => x"34010001",  2054 => x"59610004",
     2055 => x"1061000b",  2056 => x"4062000c",  2057 => x"29640028",
     2058 => x"bc411000",  2059 => x"28830018",  2060 => x"084203e8",
     2061 => x"b9600800",  2062 => x"d8600000",  2063 => x"596102d4",
     2064 => x"296102c8",  2065 => x"28210010",  2066 => x"58200064",
     2067 => x"34010001",  2068 => x"2b9d0004",  2069 => x"2b8b0008",
     2070 => x"379c0008",  2071 => x"c3a00000",  2072 => x"379cfff4",
     2073 => x"5b8b000c",  2074 => x"5b8c0008",  2075 => x"5b9d0004",
     2076 => x"78040001",  2077 => x"78050001",  2078 => x"b8606000",
     2079 => x"34020002",  2080 => x"34030002",  2081 => x"38843f18",
     2082 => x"38a55b5c",  2083 => x"b8205800",  2084 => x"fbfffa2e",
     2085 => x"29820024",  2086 => x"296102c8",  2087 => x"20430003",
     2088 => x"28210010",  2089 => x"7c640000",  2090 => x"58240038",
     2091 => x"20440008",  2092 => x"20420004",  2093 => x"7c840000",
     2094 => x"7c420000",  2095 => x"30230035",  2096 => x"58220044",
     2097 => x"58240040",  2098 => x"29610020",  2099 => x"28220010",
     2100 => x"296102c8",  2101 => x"2c210008",  2102 => x"0c41002c",
     2103 => x"2b9d0004",  2104 => x"2b8b000c",  2105 => x"2b8c0008",
     2106 => x"379c000c",  2107 => x"c3a00000",  2108 => x"379cfff8",
     2109 => x"5b8b0008",  2110 => x"5b9d0004",  2111 => x"282202c8",
     2112 => x"78040001",  2113 => x"78050001",  2114 => x"284b0010",
     2115 => x"34030002",  2116 => x"34020002",  2117 => x"38843f18",
     2118 => x"38a55c3c",  2119 => x"fbfffa0b",  2120 => x"34010000",
     2121 => x"31600005",  2122 => x"2b9d0004",  2123 => x"2b8b0008",
     2124 => x"379c0008",  2125 => x"c3a00000",  2126 => x"379cfff8",
     2127 => x"5b8b0008",  2128 => x"5b9d0004",  2129 => x"78040001",
     2130 => x"78050001",  2131 => x"b8205800",  2132 => x"34020002",
     2133 => x"34010000",  2134 => x"34030002",  2135 => x"38843f18",
     2136 => x"38a55c4c",  2137 => x"fbfff9f9",  2138 => x"29610024",
     2139 => x"44200006",  2140 => x"34020000",  2141 => x"34030001",
     2142 => x"34040002",  2143 => x"34060003",  2144 => x"e000001f",
     2145 => x"29610000",  2146 => x"29620040",  2147 => x"58220014",
     2148 => x"e000001d",  2149 => x"29650000",  2150 => x"08410374",
     2151 => x"b4a10800",  2152 => x"29650040",  2153 => x"58250014",
     2154 => x"28250368",  2155 => x"5ca30010",  2156 => x"4025001d",
     2157 => x"44a30004",  2158 => x"282102c8",  2159 => x"5ca40009",
     2160 => x"e0000005",  2161 => x"282102c8",  2162 => x"28210010",
     2163 => x"30230004",  2164 => x"e000000a",  2165 => x"28210010",
     2166 => x"30240004",  2167 => x"e0000007",  2168 => x"28210010",
     2169 => x"30260004",  2170 => x"e0000004",  2171 => x"282102c8",
     2172 => x"28210010",  2173 => x"30200004",  2174 => x"34420001",
     2175 => x"29610024",  2176 => x"4822ffe5",  2177 => x"34010000",
     2178 => x"2b9d0004",  2179 => x"2b8b0008",  2180 => x"379c0008",
     2181 => x"c3a00000",  2182 => x"379cfff4",  2183 => x"5b8b000c",
     2184 => x"5b8c0008",  2185 => x"5b9d0004",  2186 => x"282202c8",
     2187 => x"78040001",  2188 => x"78050001",  2189 => x"284b0010",
     2190 => x"34030002",  2191 => x"34020002",  2192 => x"38843f18",
     2193 => x"38a55c54",  2194 => x"b8206000",  2195 => x"fbfff9bf",
     2196 => x"41630004",  2197 => x"3401012c",  2198 => x"59610028",
     2199 => x"34020001",  2200 => x"34010bb8",  2201 => x"59610030",
     2202 => x"59600008",  2203 => x"31600035",  2204 => x"59600040",
     2205 => x"59620014",  2206 => x"20630003",  2207 => x"29610000",
     2208 => x"5c620004",  2209 => x"28230034",  2210 => x"b9800800",
     2211 => x"e0000004",  2212 => x"28230034",  2213 => x"34020000",
     2214 => x"b9800800",  2215 => x"d8600000",  2216 => x"34010000",
     2217 => x"2b9d0004",  2218 => x"2b8b000c",  2219 => x"2b8c0008",
     2220 => x"379c000c",  2221 => x"c3a00000",  2222 => x"379cfff0",
     2223 => x"5b8b0010",  2224 => x"5b8c000c",  2225 => x"5b8d0008",
     2226 => x"5b9d0004",  2227 => x"78040001",  2228 => x"78050001",
     2229 => x"2c2d0002",  2230 => x"b8205800",  2231 => x"b8406000",
     2232 => x"34010000",  2233 => x"34020002",  2234 => x"34030002",
     2235 => x"38843f18",  2236 => x"38a55ba8",  2237 => x"fbfff995",
     2238 => x"34010040",  2239 => x"4c2d0004",  2240 => x"b9600800",
     2241 => x"b9801000",  2242 => x"f8000466",  2243 => x"2b9d0004",
     2244 => x"2b8b0010",  2245 => x"2b8c000c",  2246 => x"2b8d0008",
     2247 => x"379c0010",  2248 => x"c3a00000",  2249 => x"379cfff8",
     2250 => x"5b8b0008",  2251 => x"5b9d0004",  2252 => x"78040001",
     2253 => x"78050001",  2254 => x"34020002",  2255 => x"34030002",
     2256 => x"38843f18",  2257 => x"38a55bbc",  2258 => x"b8205800",
     2259 => x"fbfff97f",  2260 => x"296102c8",  2261 => x"34020040",
     2262 => x"28210010",  2263 => x"40210004",  2264 => x"44200006",
     2265 => x"34030002",  2266 => x"44230004",  2267 => x"b9600800",
     2268 => x"f8000409",  2269 => x"3402004e",  2270 => x"b8400800",
     2271 => x"2b9d0004",  2272 => x"2b8b0008",  2273 => x"379c0008",
     2274 => x"c3a00000",  2275 => x"379cfff4",  2276 => x"5b8b000c",
     2277 => x"5b8c0008",  2278 => x"5b9d0004",  2279 => x"78040001",
     2280 => x"78050001",  2281 => x"34030002",  2282 => x"b8406000",
     2283 => x"38843f18",  2284 => x"34020002",  2285 => x"38a55bd0",
     2286 => x"b8205800",  2287 => x"fbfff963",  2288 => x"296102c8",
     2289 => x"34030000",  2290 => x"28210010",  2291 => x"28210008",
     2292 => x"44200007",  2293 => x"35630094",  2294 => x"59800008",
     2295 => x"b9600800",  2296 => x"b9801000",  2297 => x"f80005e9",
     2298 => x"34030001",  2299 => x"b8600800",  2300 => x"2b9d0004",
     2301 => x"2b8b000c",  2302 => x"2b8c0008",  2303 => x"379c000c",
     2304 => x"c3a00000",  2305 => x"379cfff8",  2306 => x"5b8b0008",
     2307 => x"5b9d0004",  2308 => x"78040001",  2309 => x"78050001",
     2310 => x"34020002",  2311 => x"34030002",  2312 => x"38843f18",
     2313 => x"38a55be4",  2314 => x"b8205800",  2315 => x"fbfff947",
     2316 => x"296102c8",  2317 => x"28220010",  2318 => x"40410004",
     2319 => x"20210002",  2320 => x"4420000b",  2321 => x"40410035",
     2322 => x"20210001",  2323 => x"44200008",  2324 => x"28410008",
     2325 => x"44200003",  2326 => x"28410040",  2327 => x"5c200004",
     2328 => x"b9600800",  2329 => x"34020009",  2330 => x"f80000a1",
     2331 => x"2b9d0004",  2332 => x"2b8b0008",  2333 => x"379c0008",
     2334 => x"c3a00000",  2335 => x"379cffdc",  2336 => x"5b8b0010",
     2337 => x"5b8c000c",  2338 => x"5b8d0008",  2339 => x"5b9d0004",
     2340 => x"28220020",  2341 => x"78040001",  2342 => x"78050001",
     2343 => x"284d0010",  2344 => x"282202c8",  2345 => x"34030002",
     2346 => x"38843f18",  2347 => x"284c0010",  2348 => x"38a55c0c",
     2349 => x"34020002",  2350 => x"b8205800",  2351 => x"fbfff923",
     2352 => x"29620318",  2353 => x"2963031c",  2354 => x"37810014",
     2355 => x"f80010df",  2356 => x"29810008",  2357 => x"5c200019",
     2358 => x"296200a0",  2359 => x"44410003",  2360 => x"296100b4",
     2361 => x"5c200008",  2362 => x"78040001",  2363 => x"b9600800",
     2364 => x"34020004",  2365 => x"34030001",  2366 => x"38843f24",
     2367 => x"fbfff913",  2368 => x"e0000013",  2369 => x"b9600800",
     2370 => x"f80011d1",  2371 => x"29a20004",  2372 => x"29810000",
     2373 => x"44400005",  2374 => x"28230034",  2375 => x"34020000",
     2376 => x"b9600800",  2377 => x"e0000004",  2378 => x"28230034",
     2379 => x"34020001",  2380 => x"b9600800",  2381 => x"d8600000",
     2382 => x"29620318",  2383 => x"b9600800",  2384 => x"f80005ac",
     2385 => x"b9600800",  2386 => x"f80005d4",  2387 => x"34010000",
     2388 => x"2b9d0004",  2389 => x"2b8b0010",  2390 => x"2b8c000c",
     2391 => x"2b8d0008",  2392 => x"379c0024",  2393 => x"c3a00000",
     2394 => x"379cfff8",  2395 => x"5b8b0008",  2396 => x"5b9d0004",
     2397 => x"78040001",  2398 => x"78050001",  2399 => x"34020002",
     2400 => x"34030002",  2401 => x"38843f18",  2402 => x"38a55c1c",
     2403 => x"b8205800",  2404 => x"fbfff8ee",  2405 => x"b9600800",
     2406 => x"f8000523",  2407 => x"34010000",  2408 => x"2b9d0004",
     2409 => x"2b8b0008",  2410 => x"379c0008",  2411 => x"c3a00000",
     2412 => x"379cffd8",  2413 => x"5b8b0010",  2414 => x"5b8c000c",
     2415 => x"5b8d0008",  2416 => x"5b9d0004",  2417 => x"78050001",
     2418 => x"b8806000",  2419 => x"78040001",  2420 => x"b8406800",
     2421 => x"34030002",  2422 => x"34020002",  2423 => x"38843f18",
     2424 => x"38a55c2c",  2425 => x"b8205800",  2426 => x"fbfff8d8",
     2427 => x"34010001",  2428 => x"45810004",  2429 => x"3401000c",
     2430 => x"5d810036",  2431 => x"e0000022",  2432 => x"296200ec",
     2433 => x"5960031c",  2434 => x"37810024",  2435 => x"4802000c",
     2436 => x"1443001f",  2437 => x"00440010",  2438 => x"3c630010",
     2439 => x"3c420010",  2440 => x"b8641800",  2441 => x"5b820028",
     2442 => x"340203e8",  2443 => x"5b830024",  2444 => x"fbfffcee",
     2445 => x"2b810028",  2446 => x"e000000d",  2447 => x"c8021000",
     2448 => x"1443001f",  2449 => x"00440010",  2450 => x"3c630010",
     2451 => x"3c420010",  2452 => x"b8641800",  2453 => x"5b820028",
     2454 => x"340203e8",  2455 => x"5b830024",  2456 => x"fbfffce2",
     2457 => x"2b810028",  2458 => x"c8010800",  2459 => x"59610318",
     2460 => x"356200e4",  2461 => x"b9600800",  2462 => x"f8001013",
     2463 => x"340c0100",  2464 => x"e0000014",  2465 => x"296102c8",
     2466 => x"b9a01000",  2467 => x"37830014",  2468 => x"28240010",
     2469 => x"b9600800",  2470 => x"340c0100",  2471 => x"3484003c",
     2472 => x"f8000416",  2473 => x"296102c8",  2474 => x"34021000",
     2475 => x"28210010",  2476 => x"2c23003c",  2477 => x"5c620007",
     2478 => x"40210004",  2479 => x"20210001",  2480 => x"44200004",
     2481 => x"b9600800",  2482 => x"34020006",  2483 => x"f8000008",
     2484 => x"b9800800",  2485 => x"2b9d0004",  2486 => x"2b8b0010",
     2487 => x"2b8c000c",  2488 => x"2b8d0008",  2489 => x"379c0028",
     2490 => x"c3a00000",  2491 => x"282302c8",  2492 => x"34040006",
     2493 => x"28630010",  2494 => x"44440004",  2495 => x"34040009",
     2496 => x"5c440008",  2497 => x"e0000004",  2498 => x"34020001",
     2499 => x"30620005",  2500 => x"e0000007",  2501 => x"34020002",
     2502 => x"30620005",  2503 => x"e0000006",  2504 => x"40630005",
     2505 => x"34020001",  2506 => x"5c620003",  2507 => x"34020066",
     2508 => x"e0000002",  2509 => x"34020064",  2510 => x"58220004",
     2511 => x"c3a00000",  2512 => x"379cfff4",  2513 => x"5b8b000c",
     2514 => x"5b8c0008",  2515 => x"5b9d0004",  2516 => x"b8205800",
     2517 => x"282102c8",  2518 => x"78050001",  2519 => x"38a53e74",
     2520 => x"282c0010",  2521 => x"34010001",  2522 => x"41820005",
     2523 => x"5c410003",  2524 => x"78050001",  2525 => x"38a5435c",
     2526 => x"78040001",  2527 => x"b9600800",  2528 => x"34020002",
     2529 => x"34030001",  2530 => x"38843f4c",  2531 => x"fbfff86f",
     2532 => x"41820005",  2533 => x"34010001",  2534 => x"5c410003",
     2535 => x"34010006",  2536 => x"e0000002",  2537 => x"34010009",
     2538 => x"59610004",  2539 => x"31800005",  2540 => x"2b9d0004",
     2541 => x"2b8b000c",  2542 => x"2b8c0008",  2543 => x"379c000c",
     2544 => x"c3a00000",  2545 => x"379cfffc",  2546 => x"5b9d0004",
     2547 => x"282202c8",  2548 => x"28420010",  2549 => x"4043002c",
     2550 => x"4460000a",  2551 => x"3463ffff",  2552 => x"78040001",
     2553 => x"3043002c",  2554 => x"38843f70",  2555 => x"34020002",
     2556 => x"34030001",  2557 => x"fbfff855",  2558 => x"34010001",
     2559 => x"e0000003",  2560 => x"fbffffd0",  2561 => x"34010000",
     2562 => x"2b9d0004",  2563 => x"379c0004",  2564 => x"c3a00000",
     2565 => x"379cffd8",  2566 => x"5b8b0018",  2567 => x"5b8c0014",
     2568 => x"5b8d0010",  2569 => x"5b8e000c",  2570 => x"5b8f0008",
     2571 => x"5b9d0004",  2572 => x"b8407000",  2573 => x"2824000c",
     2574 => x"282202c8",  2575 => x"b8205800",  2576 => x"b8607800",
     2577 => x"284d0010",  2578 => x"44800004",  2579 => x"34010003",
     2580 => x"31a1002c",  2581 => x"e000000c",  2582 => x"282202e0",
     2583 => x"44440008",  2584 => x"28220028",  2585 => x"28440018",
     2586 => x"34020000",  2587 => x"d8800000",  2588 => x"296202e0",
     2589 => x"c8220800",  2590 => x"4c20003c",  2591 => x"340c0000",
     2592 => x"e0000015",  2593 => x"29610028",  2594 => x"340203e8",
     2595 => x"28240018",  2596 => x"b9600800",  2597 => x"d8800000",
     2598 => x"596102e0",  2599 => x"296102c8",  2600 => x"29620028",
     2601 => x"4025000c",  2602 => x"1021000b",  2603 => x"28440018",
     2604 => x"bca12800",  2605 => x"b9600800",  2606 => x"08a203e8",
     2607 => x"d8800000",  2608 => x"596102d4",  2609 => x"34021000",
     2610 => x"b9600800",  2611 => x"f80003fb",  2612 => x"b8206000",
     2613 => x"45e0000e",  2614 => x"4162030d",  2615 => x"3401000c",
     2616 => x"5c41000b",  2617 => x"b9600800",  2618 => x"b9c01000",
     2619 => x"3783001c",  2620 => x"35a4003c",  2621 => x"f8000381",
     2622 => x"2da2003c",  2623 => x"34011001",  2624 => x"5c410003",
     2625 => x"34010065",  2626 => x"59610004",  2627 => x"5d800004",
     2628 => x"b9600800",  2629 => x"f8000adb",  2630 => x"e0000003",
     2631 => x"34010002",  2632 => x"59610004",  2633 => x"29620004",
     2634 => x"29610000",  2635 => x"44410002",  2636 => x"596002d4",
     2637 => x"296102c8",  2638 => x"28210010",  2639 => x"28210028",
     2640 => x"59610008",  2641 => x"b9800800",  2642 => x"2b9d0004",
     2643 => x"2b8b0018",  2644 => x"2b8c0014",  2645 => x"2b8d0010",
     2646 => x"2b8e000c",  2647 => x"2b8f0008",  2648 => x"379c0028",
     2649 => x"c3a00000",  2650 => x"b9600800",  2651 => x"34020005",
     2652 => x"f800127b",  2653 => x"b9600800",  2654 => x"596002e0",
     2655 => x"fbffff92",  2656 => x"340c0000",  2657 => x"5c20ffc0",
     2658 => x"e3ffffef",  2659 => x"379cffd8",  2660 => x"5b8b0018",
     2661 => x"5b8c0014",  2662 => x"5b8d0010",  2663 => x"5b8e000c",
     2664 => x"5b8f0008",  2665 => x"5b9d0004",  2666 => x"b8407000",
     2667 => x"2824000c",  2668 => x"282202c8",  2669 => x"b8205800",
     2670 => x"b8607800",  2671 => x"284c0010",  2672 => x"44800004",
     2673 => x"34010003",  2674 => x"3181002c",  2675 => x"e000000c",
     2676 => x"282202e0",  2677 => x"44440008",  2678 => x"28220028",
     2679 => x"28440018",  2680 => x"34020000",  2681 => x"d8800000",
     2682 => x"296202e0",  2683 => x"c8220800",  2684 => x"4c200029",
     2685 => x"340d0000",  2686 => x"e000000b",  2687 => x"34021001",
     2688 => x"b9600800",  2689 => x"f80003ad",  2690 => x"b8206800",
     2691 => x"29610028",  2692 => x"34023a98",  2693 => x"28240018",
     2694 => x"b9600800",  2695 => x"d8800000",  2696 => x"596102e0",
     2697 => x"45e0000e",  2698 => x"4162030d",  2699 => x"3401000c",
     2700 => x"5c41000b",  2701 => x"b9600800",  2702 => x"b9c01000",
     2703 => x"3783001c",  2704 => x"3584003c",  2705 => x"f800032d",
     2706 => x"2d82003c",  2707 => x"34011002",  2708 => x"5c410003",
     2709 => x"34010068",  2710 => x"59610004",  2711 => x"45a00003",
     2712 => x"34010002",  2713 => x"59610004",  2714 => x"29810028",
     2715 => x"59610008",  2716 => x"b9a00800",  2717 => x"2b9d0004",
     2718 => x"2b8b0018",  2719 => x"2b8c0014",  2720 => x"2b8d0010",
     2721 => x"2b8e000c",  2722 => x"2b8f0008",  2723 => x"379c0028",
     2724 => x"c3a00000",  2725 => x"b9600800",  2726 => x"34020005",
     2727 => x"f8001230",  2728 => x"b9600800",  2729 => x"596002e0",
     2730 => x"fbffff47",  2731 => x"340d0000",  2732 => x"5c20ffd3",
     2733 => x"e3ffffef",  2734 => x"379cfff4",  2735 => x"5b8b000c",
     2736 => x"5b8c0008",  2737 => x"5b9d0004",  2738 => x"282202c8",
     2739 => x"b8205800",  2740 => x"284c0010",  2741 => x"2822000c",
     2742 => x"44400004",  2743 => x"34010003",  2744 => x"3181002c",
     2745 => x"e000000b",  2746 => x"282302e0",  2747 => x"44620013",
     2748 => x"28220028",  2749 => x"28430018",  2750 => x"34020000",
     2751 => x"d8600000",  2752 => x"296202e0",  2753 => x"c8220800",
     2754 => x"4c200021",  2755 => x"e000000b",  2756 => x"29810000",
     2757 => x"28220000",  2758 => x"b9600800",  2759 => x"d8400000",
     2760 => x"29610028",  2761 => x"34023a98",  2762 => x"28230018",
     2763 => x"b9600800",  2764 => x"d8600000",  2765 => x"596102e0",
     2766 => x"29810000",  2767 => x"34020000",  2768 => x"28230004",
     2769 => x"b9600800",  2770 => x"d8600000",  2771 => x"34020001",
     2772 => x"5c220007",  2773 => x"34010067",  2774 => x"59610004",
     2775 => x"29810000",  2776 => x"28220008",  2777 => x"b9600800",
     2778 => x"d8400000",  2779 => x"29810028",  2780 => x"59610008",
     2781 => x"34010000",  2782 => x"2b9d0004",  2783 => x"2b8b000c",
     2784 => x"2b8c0008",  2785 => x"379c000c",  2786 => x"c3a00000",
     2787 => x"b9600800",  2788 => x"34020005",  2789 => x"f80011f2",
     2790 => x"29810000",  2791 => x"596002e0",  2792 => x"28220008",
     2793 => x"b9600800",  2794 => x"d8400000",  2795 => x"b9600800",
     2796 => x"fbffff05",  2797 => x"5c20ffd7",  2798 => x"e3ffffef",
     2799 => x"379cffd8",  2800 => x"5b8b0018",  2801 => x"5b8c0014",
     2802 => x"5b8d0010",  2803 => x"5b8e000c",  2804 => x"5b8f0008",
     2805 => x"5b9d0004",  2806 => x"b8407000",  2807 => x"2824000c",
     2808 => x"282202c8",  2809 => x"b8205800",  2810 => x"b8607800",
     2811 => x"284c0010",  2812 => x"44800004",  2813 => x"34010003",
     2814 => x"3181002c",  2815 => x"e000000c",  2816 => x"282202e0",
     2817 => x"44440008",  2818 => x"28220028",  2819 => x"28440018",
     2820 => x"34020000",  2821 => x"d8800000",  2822 => x"296202e0",
     2823 => x"c8220800",  2824 => x"4c200029",  2825 => x"340d0000",
     2826 => x"e000000b",  2827 => x"29610028",  2828 => x"29820028",
     2829 => x"28240018",  2830 => x"b9600800",  2831 => x"d8800000",
     2832 => x"596102e0",  2833 => x"34021002",  2834 => x"b9600800",
     2835 => x"f800031b",  2836 => x"b8206800",  2837 => x"45e0000e",
     2838 => x"4162030d",  2839 => x"3401000c",  2840 => x"5c41000b",
     2841 => x"b9600800",  2842 => x"b9c01000",  2843 => x"3783001c",
     2844 => x"3584003c",  2845 => x"f80002a1",  2846 => x"2d82003c",
     2847 => x"34011003",  2848 => x"5c410003",  2849 => x"3401006a",
     2850 => x"59610004",  2851 => x"45a00003",  2852 => x"34010002",
     2853 => x"59610004",  2854 => x"29810028",  2855 => x"59610008",
     2856 => x"b9a00800",  2857 => x"2b9d0004",  2858 => x"2b8b0018",
     2859 => x"2b8c0014",  2860 => x"2b8d0010",  2861 => x"2b8e000c",
     2862 => x"2b8f0008",  2863 => x"379c0028",  2864 => x"c3a00000",
     2865 => x"b9600800",  2866 => x"34020005",  2867 => x"f80011a4",
     2868 => x"b9600800",  2869 => x"596002e0",  2870 => x"fbfffebb",
     2871 => x"340d0000",  2872 => x"5c20ffd3",  2873 => x"e3ffffef",
     2874 => x"379cffec",  2875 => x"5b8b0010",  2876 => x"5b8c000c",
     2877 => x"5b8d0008",  2878 => x"5b9d0004",  2879 => x"282202c8",
     2880 => x"b8206000",  2881 => x"284b0010",  2882 => x"2822000c",
     2883 => x"44400004",  2884 => x"34010003",  2885 => x"3161002c",
     2886 => x"e000000c",  2887 => x"282302e0",  2888 => x"44620008",
     2889 => x"28220028",  2890 => x"28430018",  2891 => x"34020000",
     2892 => x"d8600000",  2893 => x"298202e0",  2894 => x"c8220800",
     2895 => x"4c2000a9",  2896 => x"340d0000",  2897 => x"e0000011",
     2898 => x"29810028",  2899 => x"29620030",  2900 => x"28230018",
     2901 => x"b9800800",  2902 => x"d8600000",  2903 => x"598102e0",
     2904 => x"34021003",  2905 => x"b9800800",  2906 => x"f80002d4",
     2907 => x"b8206800",  2908 => x"3401006c",  2909 => x"31610010",
     2910 => x"29610014",  2911 => x"44200003",  2912 => x"3401006e",
     2913 => x"31610010",  2914 => x"41660010",  2915 => x"78040001",
     2916 => x"78050001",  2917 => x"b9800800",  2918 => x"34020002",
     2919 => x"34030001",  2920 => x"38843f84",  2921 => x"38a55c80",
     2922 => x"34c6ff94",  2923 => x"fbfff6e7",  2924 => x"41620010",
     2925 => x"34010008",  2926 => x"3442ff94",  2927 => x"204200ff",
     2928 => x"5441007f",  2929 => x"78010001",  2930 => x"3c420002",
     2931 => x"38215c5c",  2932 => x"b4220800",  2933 => x"28210000",
     2934 => x"c0200000",  2935 => x"29610000",  2936 => x"34020000",
     2937 => x"34030000",  2938 => x"2825002c",  2939 => x"34040000",
     2940 => x"b9800800",  2941 => x"d8a00000",  2942 => x"5c200071",
     2943 => x"3401006d",  2944 => x"31610010",  2945 => x"29610000",
     2946 => x"34020001",  2947 => x"28230024",  2948 => x"b9800800",
     2949 => x"d8600000",  2950 => x"5c200069",  2951 => x"3401006e",
     2952 => x"31610010",  2953 => x"29610000",  2954 => x"34020001",
     2955 => x"37830014",  2956 => x"28240028",  2957 => x"b9800800",
     2958 => x"d8800000",  2959 => x"34020001",  2960 => x"5c22005f",
     2961 => x"2b810014",  2962 => x"78040001",  2963 => x"34020002",
     2964 => x"00250010",  2965 => x"3c210010",  2966 => x"5965001c",
     2967 => x"59610018",  2968 => x"34030001",  2969 => x"b9800800",
     2970 => x"38843f98",  2971 => x"fbfff6b7",  2972 => x"29650018",
     2973 => x"78040001",  2974 => x"b9800800",  2975 => x"34020002",
     2976 => x"34030001",  2977 => x"38843fbc",  2978 => x"fbfff6b0",
     2979 => x"3401006f",  2980 => x"31610010",  2981 => x"29610000",
     2982 => x"34020001",  2983 => x"28230020",  2984 => x"b9800800",
     2985 => x"d8600000",  2986 => x"5c200045",  2987 => x"34010070",
     2988 => x"31610010",  2989 => x"29610000",  2990 => x"28220030",
     2991 => x"b9800800",  2992 => x"d8400000",  2993 => x"5c20003e",
     2994 => x"34010071",  2995 => x"31610010",  2996 => x"29610000",
     2997 => x"34020002",  2998 => x"28230024",  2999 => x"b9800800",
     3000 => x"d8600000",  3001 => x"5c200036",  3002 => x"34010072",
     3003 => x"31610010",  3004 => x"29610000",  3005 => x"34020002",
     3006 => x"37830014",  3007 => x"28240028",  3008 => x"b9800800",
     3009 => x"d8800000",  3010 => x"34020001",  3011 => x"5c22002c",
     3012 => x"2b850014",  3013 => x"78040001",  3014 => x"b9800800",
     3015 => x"34020002",  3016 => x"34030001",  3017 => x"38843fe0",
     3018 => x"fbfff688",  3019 => x"2b810014",  3020 => x"78040001",
     3021 => x"34020002",  3022 => x"00250010",  3023 => x"3c210010",
     3024 => x"59650024",  3025 => x"59610020",  3026 => x"34030001",
     3027 => x"b9800800",  3028 => x"38843ff8",  3029 => x"fbfff67d",
     3030 => x"29650020",  3031 => x"78040001",  3032 => x"b9800800",
     3033 => x"34020002",  3034 => x"34030001",  3035 => x"3884401c",
     3036 => x"fbfff676",  3037 => x"34010073",  3038 => x"31610010",
     3039 => x"29610000",  3040 => x"34020002",  3041 => x"28230020",
     3042 => x"b9800800",  3043 => x"d8600000",  3044 => x"5c20000b",
     3045 => x"34010074",  3046 => x"31610010",  3047 => x"b9800800",
     3048 => x"34021004",  3049 => x"f8000245",  3050 => x"b8206800",
     3051 => x"34010069",  3052 => x"59810004",  3053 => x"34010001",
     3054 => x"59610014",  3055 => x"29610028",  3056 => x"59810008",
     3057 => x"b9a00800",  3058 => x"2b9d0004",  3059 => x"2b8b0010",
     3060 => x"2b8c000c",  3061 => x"2b8d0008",  3062 => x"379c0014",
     3063 => x"c3a00000",  3064 => x"b9800800",  3065 => x"34020005",
     3066 => x"f80010dd",  3067 => x"b9800800",  3068 => x"598002e0",
     3069 => x"fbfffdf4",  3070 => x"340d0000",  3071 => x"5c20ff53",
     3072 => x"e3fffff1",  3073 => x"379cffdc",  3074 => x"5b8b0014",
     3075 => x"5b8c0010",  3076 => x"5b8d000c",  3077 => x"5b8e0008",
     3078 => x"5b9d0004",  3079 => x"b8406800",  3080 => x"282202c8",
     3081 => x"b8205800",  3082 => x"b8607000",  3083 => x"284c0010",
     3084 => x"2822000c",  3085 => x"44400006",  3086 => x"28220028",
     3087 => x"28440018",  3088 => x"29820028",  3089 => x"d8800000",
     3090 => x"596102e0",  3091 => x"296102e0",  3092 => x"44200009",
     3093 => x"29610028",  3094 => x"34020000",  3095 => x"28240018",
     3096 => x"b9600800",  3097 => x"d8800000",  3098 => x"296202e0",
     3099 => x"c8220800",  3100 => x"4c200023",  3101 => x"45c00018",
     3102 => x"4162030d",  3103 => x"3401000c",  3104 => x"5c410015",
     3105 => x"b9600800",  3106 => x"b9a01000",  3107 => x"37830018",
     3108 => x"3584003c",  3109 => x"f8000199",  3110 => x"2d81003c",
     3111 => x"34021003",  3112 => x"5c220006",  3113 => x"41820005",
     3114 => x"34010001",  3115 => x"5c41000a",  3116 => x"3401006a",
     3117 => x"e0000007",  3118 => x"34021005",  3119 => x"5c220006",
     3120 => x"41820005",  3121 => x"34010002",  3122 => x"5c410003",
     3123 => x"3401006b",  3124 => x"59610004",  3125 => x"29810028",
     3126 => x"59610008",  3127 => x"34010000",  3128 => x"2b9d0004",
     3129 => x"2b8b0014",  3130 => x"2b8c0010",  3131 => x"2b8d000c",
     3132 => x"2b8e0008",  3133 => x"379c0024",  3134 => x"c3a00000",
     3135 => x"b9600800",  3136 => x"34020005",  3137 => x"f8001096",
     3138 => x"b9600800",  3139 => x"596002e0",  3140 => x"fbfffd8c",
     3141 => x"e3fffff2",  3142 => x"379cffd4",  3143 => x"5b8b001c",
     3144 => x"5b8c0018",  3145 => x"5b8d0014",  3146 => x"5b8e0010",
     3147 => x"5b8f000c",  3148 => x"5b900008",  3149 => x"5b9d0004",
     3150 => x"b8407000",  3151 => x"282202c8",  3152 => x"2824000c",
     3153 => x"b8205800",  3154 => x"284c0010",  3155 => x"b8607800",
     3156 => x"2d8d0048",  3157 => x"7dad0000",  3158 => x"44800004",
     3159 => x"34010003",  3160 => x"3181002c",  3161 => x"e0000012",
     3162 => x"282202e0",  3163 => x"44440022",  3164 => x"28220028",
     3165 => x"28440018",  3166 => x"34020000",  3167 => x"d8800000",
     3168 => x"296202e0",  3169 => x"c8220800",  3170 => x"4c20003f",
     3171 => x"e000001a",  3172 => x"29810000",  3173 => x"28240030",
     3174 => x"b9600800",  3175 => x"d8800000",  3176 => x"b9600800",
     3177 => x"fbfffd88",  3178 => x"4420002d",  3179 => x"45a00008",
     3180 => x"29810000",  3181 => x"34020000",  3182 => x"34030000",
     3183 => x"2825002c",  3184 => x"34040000",  3185 => x"b9600800",
     3186 => x"d8a00000",  3187 => x"2981004c",  3188 => x"29700028",
     3189 => x"340203e8",  3190 => x"f8003eec",  3191 => x"2a050018",
     3192 => x"b8202000",  3193 => x"b8801000",  3194 => x"b9600800",
     3195 => x"d8a00000",  3196 => x"596102e0",  3197 => x"45e00018",
     3198 => x"4162030d",  3199 => x"3401000c",  3200 => x"5c410015",
     3201 => x"b9600800",  3202 => x"b9c01000",  3203 => x"37830020",
     3204 => x"3584003c",  3205 => x"f8000139",  3206 => x"2d82003c",
     3207 => x"34011004",  3208 => x"5c41000d",  3209 => x"45a00005",
     3210 => x"29810000",  3211 => x"28220030",  3212 => x"b9600800",
     3213 => x"d8400000",  3214 => x"41820005",  3215 => x"34010001",
     3216 => x"5c410003",  3217 => x"3401006b",  3218 => x"e0000002",
     3219 => x"34010068",  3220 => x"59610004",  3221 => x"29810028",
     3222 => x"59610008",  3223 => x"34010000",  3224 => x"2b9d0004",
     3225 => x"2b8b001c",  3226 => x"2b8c0018",  3227 => x"2b8d0014",
     3228 => x"2b8e0010",  3229 => x"2b8f000c",  3230 => x"2b900008",
     3231 => x"379c002c",  3232 => x"c3a00000",  3233 => x"b9600800",
     3234 => x"34020005",  3235 => x"f8001034",  3236 => x"596002e0",
     3237 => x"45a0ffc3",  3238 => x"e3ffffbe",  3239 => x"379cfff0",
     3240 => x"5b8b0010",  3241 => x"5b8c000c",  3242 => x"5b8d0008",
     3243 => x"5b9d0004",  3244 => x"282202c8",  3245 => x"340d0001",
     3246 => x"b8206000",  3247 => x"284b0010",  3248 => x"29620000",
     3249 => x"596d0008",  3250 => x"2842000c",  3251 => x"d8400000",
     3252 => x"41610005",  3253 => x"34020000",  3254 => x"5c2d0005",
     3255 => x"34021005",  3256 => x"b9800800",  3257 => x"f8000175",
     3258 => x"b8201000",  3259 => x"34010001",  3260 => x"59610040",
     3261 => x"3401ffff",  3262 => x"5c400009",  3263 => x"41620005",
     3264 => x"34010002",  3265 => x"5c410003",  3266 => x"34010009",
     3267 => x"e0000002",  3268 => x"34010006",  3269 => x"59810004",
     3270 => x"34010000",  3271 => x"2b9d0004",  3272 => x"2b8b0010",
     3273 => x"2b8c000c",  3274 => x"2b8d0008",  3275 => x"379c0010",
     3276 => x"c3a00000",  3277 => x"00430018",  3278 => x"30220003",
     3279 => x"30230000",  3280 => x"00430010",  3281 => x"30230001",
     3282 => x"00430008",  3283 => x"30230002",  3284 => x"c3a00000",
     3285 => x"40220000",  3286 => x"40230003",  3287 => x"3c420018",
     3288 => x"b8621000",  3289 => x"40230001",  3290 => x"40210002",
     3291 => x"3c630010",  3292 => x"3c210008",  3293 => x"b8431000",
     3294 => x"b8410800",  3295 => x"c3a00000",  3296 => x"40220000",
     3297 => x"40210001",  3298 => x"3c420008",  3299 => x"b8410800",
     3300 => x"c3a00000",  3301 => x"379cfff0",  3302 => x"5b8b0010",
     3303 => x"5b8c000c",  3304 => x"5b8d0008",  3305 => x"5b9d0004",
     3306 => x"28230020",  3307 => x"282202c8",  3308 => x"b8205800",
     3309 => x"2863000c",  3310 => x"28420010",  3311 => x"282c003c",
     3312 => x"4064000e",  3313 => x"340300ba",  3314 => x"48830018",
     3315 => x"28420000",  3316 => x"28430004",  3317 => x"34020001",
     3318 => x"d8600000",  3319 => x"ec016800",  3320 => x"b9600800",
     3321 => x"f8000994",  3322 => x"29610020",  3323 => x"c80d6800",
     3324 => x"21ad002e",  3325 => x"2821000c",  3326 => x"35ad0006",
     3327 => x"4021000e",  3328 => x"45a1000a",  3329 => x"78010001",
     3330 => x"b9a01000",  3331 => x"38214040",  3332 => x"f80024eb",
     3333 => x"29610020",  3334 => x"21ad00ff",  3335 => x"2821000c",
     3336 => x"302d000e",  3337 => x"318d0030",  3338 => x"3401004e",
     3339 => x"0d810002",  3340 => x"34010003",  3341 => x"0d810040",
     3342 => x"3401000a",  3343 => x"0d810042",  3344 => x"34010800",
     3345 => x"0d810044",  3346 => x"340130de",  3347 => x"0d810046",
     3348 => x"3401ad01",  3349 => x"0d810048",  3350 => x"34012000",
     3351 => x"0d81004a",  3352 => x"296102c8",  3353 => x"28220010",
     3354 => x"28430014",  3355 => x"40410004",  3356 => x"44600002",
     3357 => x"38210004",  3358 => x"28420008",  3359 => x"44400002",
     3360 => x"38210008",  3361 => x"0d81004c",  3362 => x"2b9d0004",
     3363 => x"2b8b0010",  3364 => x"2b8c000c",  3365 => x"2b8d0008",
     3366 => x"379c0010",  3367 => x"c3a00000",  3368 => x"379cfff4",
     3369 => x"5b8b000c",  3370 => x"5b8c0008",  3371 => x"5b9d0004",
     3372 => x"b8205800",  3373 => x"34210040",  3374 => x"b8406000",
     3375 => x"fbffffb1",  3376 => x"2d650044",  3377 => x"2d640046",
     3378 => x"78070001",  3379 => x"3ca50008",  3380 => x"00860008",
     3381 => x"38e75a34",  3382 => x"b8a62800",  3383 => x"28e60000",
     3384 => x"64210003",  3385 => x"2d630048",  3386 => x"e4a62800",
     3387 => x"2d62004a",  3388 => x"a0250800",  3389 => x"44200010",
     3390 => x"3c840008",  3391 => x"00610008",  3392 => x"2084ffff",
     3393 => x"b8812000",  3394 => x"206300ff",  3395 => x"3801dead",
     3396 => x"e4812000",  3397 => x"64630001",  3398 => x"a0831800",
     3399 => x"44600006",  3400 => x"34012000",  3401 => x"5c410004",
     3402 => x"3561004c",  3403 => x"fbffff95",  3404 => x"59810024",
     3405 => x"2b9d0004",  3406 => x"2b8b000c",  3407 => x"2b8c0008",
     3408 => x"379c000c",  3409 => x"c3a00000",  3410 => x"379cfff0",
     3411 => x"5b8b0010",  3412 => x"5b8c000c",  3413 => x"5b8d0008",
     3414 => x"5b9d0004",  3415 => x"b8206000",  3416 => x"282102c8",
     3417 => x"204dffff",  3418 => x"28210010",  3419 => x"40250005",
     3420 => x"44a00003",  3421 => x"34012000",  3422 => x"5da1000a",
     3423 => x"78040001",  3424 => x"b9800800",  3425 => x"34020005",
     3426 => x"34030001",  3427 => x"38844058",  3428 => x"b9a03000",
     3429 => x"fbfff4ed",  3430 => x"34010000",  3431 => x"e0000051",
     3432 => x"298b003c",  3433 => x"34030008",  3434 => x"41610000",
     3435 => x"202100f0",  3436 => x"3821000c",  3437 => x"31610000",
     3438 => x"34010005",  3439 => x"31610020",  3440 => x"29820020",
     3441 => x"35610022",  3442 => x"28420014",  3443 => x"f8003e50",
     3444 => x"29810020",  3445 => x"28210014",  3446 => x"2c210008",
     3447 => x"0d6d0036",  3448 => x"00220008",  3449 => x"3161002b",
     3450 => x"34010003",  3451 => x"0d61002c",  3452 => x"34010800",
     3453 => x"0d610030",  3454 => x"340130de",  3455 => x"0d610032",
     3456 => x"3401ad01",  3457 => x"0d610034",  3458 => x"3162002a",
     3459 => x"34011003",  3460 => x"45a10005",  3461 => x"34011004",
     3462 => x"34020008",  3463 => x"5da1002d",  3464 => x"e0000017",
     3465 => x"298102c8",  3466 => x"35620038",  3467 => x"28210010",
     3468 => x"28230014",  3469 => x"44600005",  3470 => x"40210034",
     3471 => x"31610038",  3472 => x"30400001",  3473 => x"e0000007",
     3474 => x"40210034",  3475 => x"3c210008",  3476 => x"38210001",
     3477 => x"00230008",  3478 => x"31630038",  3479 => x"30410001",
     3480 => x"298102c8",  3481 => x"28220010",  3482 => x"3561003a",
     3483 => x"28420030",  3484 => x"fbffff31",  3485 => x"34020014",
     3486 => x"e0000016",  3487 => x"298102c8",  3488 => x"28220010",
     3489 => x"35610038",  3490 => x"2842001c",  3491 => x"fbffff2a",
     3492 => x"298102c8",  3493 => x"28220010",  3494 => x"3561003c",
     3495 => x"28420018",  3496 => x"fbffff25",  3497 => x"298102c8",
     3498 => x"28220010",  3499 => x"35610040",  3500 => x"28420024",
     3501 => x"fbffff20",  3502 => x"298102c8",  3503 => x"28220010",
     3504 => x"35610044",  3505 => x"28420020",  3506 => x"fbffff1b",
     3507 => x"34020018",  3508 => x"34410030",  3509 => x"31600002",
     3510 => x"31610003",  3511 => x"0d62002e",  3512 => x"2b9d0004",
     3513 => x"2b8b0010",  3514 => x"2b8c000c",  3515 => x"2b8d0008",
     3516 => x"379c0010",  3517 => x"c3a00000",  3518 => x"379cffec",
     3519 => x"5b8b0014",  3520 => x"5b8c0010",  3521 => x"5b8d000c",
     3522 => x"5b8e0008",  3523 => x"5b9d0004",  3524 => x"b8405800",
     3525 => x"b8607000",  3526 => x"34420022",  3527 => x"b8206000",
     3528 => x"b8600800",  3529 => x"34030008",  3530 => x"b8806800",
     3531 => x"f8003df8",  3532 => x"3561002a",  3533 => x"fbffff13",
     3534 => x"0dc10008",  3535 => x"3561002c",  3536 => x"fbffff10",
     3537 => x"b8202800",  3538 => x"34040003",  3539 => x"2d630030",
     3540 => x"2d620032",  3541 => x"2d610034",  3542 => x"44a40007",
     3543 => x"78040001",  3544 => x"b9800800",  3545 => x"34020005",
     3546 => x"34030001",  3547 => x"3884408c",  3548 => x"e0000022",
     3549 => x"3c650008",  3550 => x"78040001",  3551 => x"00430008",
     3552 => x"38845a34",  3553 => x"b8a32800",  3554 => x"28830000",
     3555 => x"44a30007",  3556 => x"78040001",  3557 => x"b9800800",
     3558 => x"34020005",  3559 => x"34030001",  3560 => x"388440dc",
     3561 => x"e0000015",  3562 => x"3c450008",  3563 => x"00230008",
     3564 => x"20a5ffff",  3565 => x"b8a32800",  3566 => x"3802dead",
     3567 => x"44a20007",  3568 => x"78040001",  3569 => x"b9800800",
     3570 => x"34020005",  3571 => x"34030001",  3572 => x"38844114",
     3573 => x"e0000009",  3574 => x"202500ff",  3575 => x"34010001",
     3576 => x"44a10008",  3577 => x"78040001",  3578 => x"b9800800",
     3579 => x"34020005",  3580 => x"34030001",  3581 => x"38844158",
     3582 => x"fbfff454",  3583 => x"e0000028",  3584 => x"2d610036",
     3585 => x"45a00002",  3586 => x"0da10000",  3587 => x"34021003",
     3588 => x"44220004",  3589 => x"34021004",  3590 => x"5c220021",
     3591 => x"e0000012",  3592 => x"298102c8",  3593 => x"356e0038",
     3594 => x"282d0010",  3595 => x"b9c00800",  3596 => x"fbfffed4",
     3597 => x"202100ff",  3598 => x"0da10048",  3599 => x"b9c00800",
     3600 => x"fbfffed0",  3601 => x"00210008",  3602 => x"31a10050",
     3603 => x"3561003a",  3604 => x"fbfffec1",  3605 => x"298202c8",
     3606 => x"28420010",  3607 => x"5841004c",  3608 => x"e000000f",
     3609 => x"298102c8",  3610 => x"282c0010",  3611 => x"35610038",
     3612 => x"fbfffeb9",  3613 => x"59810058",  3614 => x"3561003c",
     3615 => x"fbfffeb6",  3616 => x"59810054",  3617 => x"35610040",
     3618 => x"fbfffeb3",  3619 => x"59810060",  3620 => x"35610044",
     3621 => x"fbfffeb0",  3622 => x"5981005c",  3623 => x"2b9d0004",
     3624 => x"2b8b0014",  3625 => x"2b8c0010",  3626 => x"2b8d000c",
     3627 => x"2b8e0008",  3628 => x"379c0014",  3629 => x"c3a00000",
     3630 => x"379cfff4",  3631 => x"5b8b000c",  3632 => x"5b8c0008",
     3633 => x"5b9d0004",  3634 => x"2042ffff",  3635 => x"b8205800",
     3636 => x"fbffff1e",  3637 => x"b8206000",  3638 => x"29610024",
     3639 => x"29630070",  3640 => x"29620034",  3641 => x"2827000c",
     3642 => x"b5831800",  3643 => x"b9600800",  3644 => x"356400f8",
     3645 => x"34050000",  3646 => x"34060000",  3647 => x"d8e00000",
     3648 => x"78080001",  3649 => x"390867c4",  3650 => x"4c2c000b",
     3651 => x"29050030",  3652 => x"78040001",  3653 => x"b9600800",
     3654 => x"34020005",  3655 => x"34030001",  3656 => x"3884419c",
     3657 => x"3406000c",  3658 => x"fbfff408",  3659 => x"3401ffff",
     3660 => x"e000000f",  3661 => x"296600f8",  3662 => x"296700fc",
     3663 => x"29080030",  3664 => x"78040001",  3665 => x"b9600800",
     3666 => x"34020005",  3667 => x"34030001",  3668 => x"388441bc",
     3669 => x"b9802800",  3670 => x"fbfff3fc",  3671 => x"2961036c",
     3672 => x"34210001",  3673 => x"5961036c",  3674 => x"34010000",
     3675 => x"2b9d0004",  3676 => x"2b8b000c",  3677 => x"2b8c0008",
     3678 => x"379c000c",  3679 => x"c3a00000",  3680 => x"78020001",
     3681 => x"384267c0",  3682 => x"58410000",  3683 => x"c3a00000",
     3684 => x"379cffe8",  3685 => x"5b8b0018",  3686 => x"5b8c0014",
     3687 => x"5b8d0010",  3688 => x"5b8e000c",  3689 => x"5b8f0008",
     3690 => x"5b9d0004",  3691 => x"282b0014",  3692 => x"b8206800",
     3693 => x"45600014",  3694 => x"780c0001",  3695 => x"398c92a4",
     3696 => x"29810000",  3697 => x"34020001",  3698 => x"f8001229",
     3699 => x"34020000",  3700 => x"31a0001c",  3701 => x"b9600800",
     3702 => x"34030110",  3703 => x"296f00f0",  3704 => x"296e00f4",
     3705 => x"296d00f8",  3706 => x"f8003dc7",  3707 => x"29810000",
     3708 => x"596f00f0",  3709 => x"596e00f4",  3710 => x"596d00f8",
     3711 => x"34020000",  3712 => x"f800121b",  3713 => x"2b9d0004",
     3714 => x"2b8b0018",  3715 => x"2b8c0014",  3716 => x"2b8d0010",
     3717 => x"2b8e000c",  3718 => x"2b8f0008",  3719 => x"379c0018",
     3720 => x"c3a00000",  3721 => x"379cffec",  3722 => x"5b8b0014",
     3723 => x"5b8c0010",  3724 => x"5b8d000c",  3725 => x"5b8e0008",
     3726 => x"5b9d0004",  3727 => x"b8206800",  3728 => x"282102c8",
     3729 => x"780e0001",  3730 => x"39ce92a4",  3731 => x"282c0010",
     3732 => x"29c10000",  3733 => x"34020001",  3734 => x"29ab0014",
     3735 => x"f8001204",  3736 => x"29810000",  3737 => x"34020000",
     3738 => x"34030000",  3739 => x"2826001c",  3740 => x"35640028",
     3741 => x"b9a00800",  3742 => x"3565002c",  3743 => x"d8c00000",
     3744 => x"3402ffff",  3745 => x"5c200039",  3746 => x"29810000",
     3747 => x"34020000",  3748 => x"28230034",  3749 => x"b9a00800",
     3750 => x"d8600000",  3751 => x"34030010",  3752 => x"35a20358",
     3753 => x"b9600800",  3754 => x"f8003ec9",  3755 => x"29810000",
     3756 => x"596000a8",  3757 => x"28220018",  3758 => x"34010000",
     3759 => x"d8400000",  3760 => x"34010002",  3761 => x"59610014",
     3762 => x"29810058",  3763 => x"2d820054",  3764 => x"59600088",
     3765 => x"3c210010",  3766 => x"b8220800",  3767 => x"59610018",
     3768 => x"29810060",  3769 => x"2d82005c",  3770 => x"3c210010",
     3771 => x"b8220800",  3772 => x"5961001c",  3773 => x"2981001c",
     3774 => x"2d820018",  3775 => x"3c210010",  3776 => x"b8220800",
     3777 => x"59610020",  3778 => x"29810024",  3779 => x"2d820020",
     3780 => x"3c210010",  3781 => x"b8220800",  3782 => x"78020001",
     3783 => x"59610024",  3784 => x"384241e0",  3785 => x"356100c0",
     3786 => x"f8003e09",  3787 => x"29610010",  3788 => x"34020000",
     3789 => x"596000b8",  3790 => x"38210001",  3791 => x"59610010",
     3792 => x"78010001",  3793 => x"382167c0",  3794 => x"28210000",
     3795 => x"596100bc",  3796 => x"78010001",  3797 => x"38217a80",
     3798 => x"58200000",  3799 => x"29c10000",  3800 => x"f80011c3",
     3801 => x"34020000",  3802 => x"b8400800",  3803 => x"2b9d0004",
     3804 => x"2b8b0014",  3805 => x"2b8c0010",  3806 => x"2b8d000c",
     3807 => x"2b8e0008",  3808 => x"379c0014",  3809 => x"c3a00000",
     3810 => x"28460000",  3811 => x"28450004",  3812 => x"28440008",
     3813 => x"28210014",  3814 => x"28420010",  3815 => x"58260030",
     3816 => x"58220040",  3817 => x"34020001",  3818 => x"58250034",
     3819 => x"58240038",  3820 => x"5822003c",  3821 => x"28670000",
     3822 => x"28660004",  3823 => x"28650008",  3824 => x"2864000c",
     3825 => x"28630010",  3826 => x"58270044",  3827 => x"58260048",
     3828 => x"5825004c",  3829 => x"58240050",  3830 => x"58230054",
     3831 => x"78010001",  3832 => x"38217a80",  3833 => x"58220000",
     3834 => x"34010000",  3835 => x"c3a00000",  3836 => x"379cfff8",
     3837 => x"5b8b0008",  3838 => x"5b9d0004",  3839 => x"282500b0",
     3840 => x"282400b4",  3841 => x"282300b8",  3842 => x"282b0014",
     3843 => x"282700a8",  3844 => x"282600ac",  3845 => x"59650060",
     3846 => x"59640064",  3847 => x"282500bc",  3848 => x"282400c0",
     3849 => x"59630068",  3850 => x"282300c4",  3851 => x"282100cc",
     3852 => x"59670058",  3853 => x"59640070",  3854 => x"5961007c",
     3855 => x"34010001",  3856 => x"59610078",  3857 => x"1441001f",
     3858 => x"59630074",  3859 => x"5966005c",  3860 => x"5965006c",
     3861 => x"34030000",  3862 => x"340403e8",  3863 => x"f8003bd7",
     3864 => x"1423001f",  3865 => x"2063ffff",  3866 => x"b4621000",
     3867 => x"f4621800",  3868 => x"00420010",  3869 => x"b4610800",
     3870 => x"3c210010",  3871 => x"b8221000",  3872 => x"34010000",
     3873 => x"59620074",  3874 => x"2b9d0004",  3875 => x"2b8b0008",
     3876 => x"379c0008",  3877 => x"c3a00000",  3878 => x"379cffbc",
     3879 => x"5b8b003c",  3880 => x"5b8c0038",  3881 => x"5b8d0034",
     3882 => x"5b8e0030",  3883 => x"5b8f002c",  3884 => x"5b900028",
     3885 => x"5b910024",  3886 => x"5b920020",  3887 => x"5b93001c",
     3888 => x"5b940018",  3889 => x"5b950014",  3890 => x"5b960010",
     3891 => x"5b97000c",  3892 => x"5b980008",  3893 => x"5b9d0004",
     3894 => x"b8206000",  3895 => x"282102c8",  3896 => x"298b0014",
     3897 => x"282e0010",  3898 => x"78010001",  3899 => x"38217a80",
     3900 => x"28210000",  3901 => x"44200283",  3902 => x"2963003c",
     3903 => x"44600007",  3904 => x"29610050",  3905 => x"44200005",
     3906 => x"29610064",  3907 => x"44200003",  3908 => x"29610078",
     3909 => x"5c200011",  3910 => x"78010001",  3911 => x"38217a84",
     3912 => x"28220000",  3913 => x"34420001",  3914 => x"58220000",
     3915 => x"34010005",  3916 => x"4c220274",  3917 => x"29640050",
     3918 => x"29650064",  3919 => x"29660078",  3920 => x"78010001",
     3921 => x"78020001",  3922 => x"38425cbc",  3923 => x"38214200",
     3924 => x"f800229b",  3925 => x"e000026b",  3926 => x"29c10000",
     3927 => x"28230038",  3928 => x"44600004",  3929 => x"b9600800",
     3930 => x"34020000",  3931 => x"d8600000",  3932 => x"78010001",
     3933 => x"382192a4",  3934 => x"28210000",  3935 => x"34020001",
     3936 => x"f800113b",  3937 => x"78010001",  3938 => x"38217a84",
     3939 => x"58200000",  3940 => x"296100b8",  3941 => x"356200fc",
     3942 => x"34210001",  3943 => x"596100b8",  3944 => x"29810028",
     3945 => x"28230000",  3946 => x"b9800800",  3947 => x"d8600000",
     3948 => x"78010001",  3949 => x"38217a80",  3950 => x"58200000",
     3951 => x"29660030",  3952 => x"29670034",  3953 => x"29680038",
     3954 => x"2965006c",  3955 => x"29640074",  3956 => x"29610070",
     3957 => x"c8a62800",  3958 => x"c8882000",  3959 => x"c8270800",
     3960 => x"e0000002",  3961 => x"348403e8",  3962 => x"b8201800",
     3963 => x"3421ffff",  3964 => x"4804fffd",  3965 => x"b8a00800",
     3966 => x"78050001",  3967 => x"38a55a2c",  3968 => x"28a20000",
     3969 => x"e0000002",  3970 => x"b4621800",  3971 => x"b8205000",
     3972 => x"3421ffff",  3973 => x"4803fffd",  3974 => x"29610044",
     3975 => x"29650058",  3976 => x"29620060",  3977 => x"2969005c",
     3978 => x"c8a12800",  3979 => x"2961004c",  3980 => x"c8410800",
     3981 => x"29620048",  3982 => x"c9224800",  3983 => x"e0000002",
     3984 => x"342103e8",  3985 => x"b9201000",  3986 => x"3529ffff",
     3987 => x"4801fffd",  3988 => x"78090001",  3989 => x"39295a2c",
     3990 => x"292d0000",  3991 => x"e0000002",  3992 => x"b44d1000",
     3993 => x"b8a04800",  3994 => x"34a5ffff",  3995 => x"4802fffd",
     3996 => x"c8810800",  3997 => x"c9495000",  3998 => x"c8622000",
     3999 => x"e0000002",  4000 => x"342103e8",  4001 => x"b8801000",
     4002 => x"3484ffff",  4003 => x"4801fffd",  4004 => x"78040001",
     4005 => x"38845a2c",  4006 => x"b9401800",  4007 => x"28850000",
     4008 => x"e0000002",  4009 => x"b4451000",  4010 => x"b8602000",
     4011 => x"3463ffff",  4012 => x"4802fffd",  4013 => x"59610094",
     4014 => x"78010001",  4015 => x"3821758c",  4016 => x"59620090",
     4017 => x"28210000",  4018 => x"29820018",  4019 => x"5964008c",
     4020 => x"b8220800",  4021 => x"00210010",  4022 => x"2021000f",
     4023 => x"44200032",  4024 => x"780d0001",  4025 => x"39ad4230",
     4026 => x"78050001",  4027 => x"b9800800",  4028 => x"34020004",
     4029 => x"34030002",  4030 => x"b9a02000",  4031 => x"38a54240",
     4032 => x"fbfff292",  4033 => x"29660044",  4034 => x"29670048",
     4035 => x"2968004c",  4036 => x"78050001",  4037 => x"b9800800",
     4038 => x"34020004",  4039 => x"34030002",  4040 => x"b9a02000",
     4041 => x"38a5424c",  4042 => x"fbfff288",  4043 => x"29660058",
     4044 => x"2967005c",  4045 => x"29680060",  4046 => x"78050001",
     4047 => x"b9800800",  4048 => x"34020004",  4049 => x"34030002",
     4050 => x"b9a02000",  4051 => x"38a54258",  4052 => x"fbfff27e",
     4053 => x"2966006c",  4054 => x"29670070",  4055 => x"29680074",
     4056 => x"78050001",  4057 => x"b9800800",  4058 => x"34020004",
     4059 => x"34030002",  4060 => x"b9a02000",  4061 => x"38a54264",
     4062 => x"fbfff274",  4063 => x"2966008c",  4064 => x"29670090",
     4065 => x"29680094",  4066 => x"78050001",  4067 => x"b9800800",
     4068 => x"34020004",  4069 => x"34030002",  4070 => x"b9a02000",
     4071 => x"38a54270",  4072 => x"fbfff26a",  4073 => x"2962008c",
     4074 => x"78050001",  4075 => x"38a55a38",  4076 => x"28a40000",
     4077 => x"1441001f",  4078 => x"340300e8",  4079 => x"f8003aff",
     4080 => x"b8406800",  4081 => x"29620090",  4082 => x"b8207800",
     4083 => x"34030000",  4084 => x"1441001f",  4085 => x"340403e8",
     4086 => x"f8003af8",  4087 => x"29660094",  4088 => x"b5a21800",
     4089 => x"f5a36800",  4090 => x"14c2001f",  4091 => x"b5e10800",
     4092 => x"b4663000",  4093 => x"b5a10800",  4094 => x"f4661800",
     4095 => x"b4220800",  4096 => x"29650018",  4097 => x"29620020",
     4098 => x"2964001c",  4099 => x"b4610800",  4100 => x"29630024",
     4101 => x"b4a21000",  4102 => x"b4441000",  4103 => x"b4431000",
     4104 => x"1444001f",  4105 => x"297600a0",  4106 => x"297400a4",
     4107 => x"596100a0",  4108 => x"596600a4",  4109 => x"48810004",
     4110 => x"5c810005",  4111 => x"54460002",  4112 => x"e0000003",
     4113 => x"596400a0",  4114 => x"596200a4",  4115 => x"296600a4",
     4116 => x"296100a0",  4117 => x"1477001f",  4118 => x"c8c21000",
     4119 => x"f4463000",  4120 => x"c8240800",  4121 => x"c8260800",
     4122 => x"b4652000",  4123 => x"14a6001f",  4124 => x"f4641800",
     4125 => x"b6e6b800",  4126 => x"b477b800",  4127 => x"004d0001",
     4128 => x"3c23001f",  4129 => x"00250001",  4130 => x"b86d6800",
     4131 => x"b48d6800",  4132 => x"f48d2000",  4133 => x"b6e5b800",
     4134 => x"b497b800",  4135 => x"29640028",  4136 => x"1483001f",
     4137 => x"f8003ac5",  4138 => x"14350008",  4139 => x"1421001f",
     4140 => x"b5b5a800",  4141 => x"f5b56800",  4142 => x"b6e10800",
     4143 => x"b5a1b800",  4144 => x"29620030",  4145 => x"29610044",
     4146 => x"29720038",  4147 => x"29630034",  4148 => x"c8411000",
     4149 => x"2961004c",  4150 => x"ca419000",  4151 => x"29610048",
     4152 => x"c8611800",  4153 => x"e0000002",  4154 => x"365203e8",
     4155 => x"b8606800",  4156 => x"3463ffff",  4157 => x"4812fffd",
     4158 => x"78090001",  4159 => x"39295a2c",  4160 => x"29210000",
     4161 => x"e0000002",  4162 => x"b5a16800",  4163 => x"b8408800",
     4164 => x"3442ffff",  4165 => x"480dfffd",  4166 => x"378f0040",
     4167 => x"340203e8",  4168 => x"b9e00800",  4169 => x"5b970040",
     4170 => x"5b950044",  4171 => x"fbfff62f",  4172 => x"78030001",
     4173 => x"38635a2c",  4174 => x"28620000",  4175 => x"b8208000",
     4176 => x"b9e00800",  4177 => x"fbfff629",  4178 => x"2b820044",
     4179 => x"b42d6800",  4180 => x"b6509000",  4181 => x"b6221000",
     4182 => x"340103e7",  4183 => x"e0000002",  4184 => x"3652fc18",
     4185 => x"b9a08800",  4186 => x"ba408000",  4187 => x"35ad0001",
     4188 => x"4a41fffc",  4189 => x"78040001",  4190 => x"78050001",
     4191 => x"38845a3c",  4192 => x"38a55a40",  4193 => x"b8400800",
     4194 => x"28830000",  4195 => x"28a20000",  4196 => x"e0000002",
     4197 => x"b6228800",  4198 => x"b8207800",  4199 => x"ba206800",
     4200 => x"34210001",  4201 => x"4a23fffc",  4202 => x"2961002c",
     4203 => x"340203e8",  4204 => x"b9e0c000",  4205 => x"342103e7",
     4206 => x"f8003aa7",  4207 => x"b8209800",  4208 => x"4c110008",
     4209 => x"ba200800",  4210 => x"ba601000",  4211 => x"f8003acf",
     4212 => x"4420000a",  4213 => x"083003e8",  4214 => x"ca216800",
     4215 => x"b6128000",  4216 => x"4da00006",  4217 => x"78090001",
     4218 => x"39295a2c",  4219 => x"29210000",  4220 => x"35efffff",
     4221 => x"b5a16800",  4222 => x"3401ffff",  4223 => x"5de10007",
     4224 => x"4c0d0006",  4225 => x"78020001",  4226 => x"38425a40",
     4227 => x"28410000",  4228 => x"340f0000",  4229 => x"b5a16800",
     4230 => x"4da00007",  4231 => x"c8130800",  4232 => x"482d0005",
     4233 => x"5de00004",  4234 => x"b5b36800",  4235 => x"0a73fc18",
     4236 => x"b6138000",  4237 => x"78050001",  4238 => x"38a55a38",
     4239 => x"28a40000",  4240 => x"1701001f",  4241 => x"bb001000",
     4242 => x"340300e8",  4243 => x"f8003a5b",  4244 => x"b820c000",
     4245 => x"1621001f",  4246 => x"b8409800",  4247 => x"34030000",
     4248 => x"340403e8",  4249 => x"ba201000",  4250 => x"f8003a54",
     4251 => x"b6621800",  4252 => x"f6639800",  4253 => x"1642001f",
     4254 => x"b7010800",  4255 => x"b4729000",  4256 => x"b6610800",
     4257 => x"b4220800",  4258 => x"f4721800",  4259 => x"78020001",
     4260 => x"384267c0",  4261 => x"b4611800",  4262 => x"28410000",
     4263 => x"596300e8",  4264 => x"34020000",  4265 => x"596100bc",
     4266 => x"29c10000",  4267 => x"597200ec",  4268 => x"597700b0",
     4269 => x"28230004",  4270 => x"597500b4",  4271 => x"b9800800",
     4272 => x"d8600000",  4273 => x"34020001",  4274 => x"4422000c",
     4275 => x"78040001",  4276 => x"b9800800",  4277 => x"34020004",
     4278 => x"34030001",  4279 => x"3884427c",  4280 => x"fbfff19a",
     4281 => x"29c10000",  4282 => x"34020000",  4283 => x"28230034",
     4284 => x"b9800800",  4285 => x"d8600000",  4286 => x"29c10000",
     4287 => x"28210010",  4288 => x"d8200000",  4289 => x"5c200007",
     4290 => x"29630010",  4291 => x"3402fffd",  4292 => x"a0621000",
     4293 => x"59620010",  4294 => x"5de10009",  4295 => x"e000000a",
     4296 => x"78040001",  4297 => x"b9800800",  4298 => x"34020004",
     4299 => x"34030001",  4300 => x"388442a0",  4301 => x"fbfff185",
     4302 => x"e00000e7",  4303 => x"34010002",  4304 => x"e0000003",
     4305 => x"45af0003",  4306 => x"34010001",  4307 => x"59610014",
     4308 => x"78040001",  4309 => x"b9800800",  4310 => x"34020004",
     4311 => x"b9e02800",  4312 => x"b9a03000",  4313 => x"34030002",
     4314 => x"388442ac",  4315 => x"ba003800",  4316 => x"fbfff176",
     4317 => x"29620014",  4318 => x"78010001",  4319 => x"38215ca4",
     4320 => x"3c420002",  4321 => x"78060001",  4322 => x"b4220800",
     4323 => x"28250000",  4324 => x"29610010",  4325 => x"38c65a24",
     4326 => x"20210002",  4327 => x"44200003",  4328 => x"78060001",
     4329 => x"38c641f0",  4330 => x"78040001",  4331 => x"b9800800",
     4332 => x"34020004",  4333 => x"34030001",  4334 => x"388442cc",
     4335 => x"fbfff163",  4336 => x"29620014",  4337 => x"78010001",
     4338 => x"38215ca4",  4339 => x"3c420002",  4340 => x"b4221000",
     4341 => x"28420000",  4342 => x"356100c0",  4343 => x"f8003bdc",
     4344 => x"29620014",  4345 => x"34010004",  4346 => x"3442ffff",
     4347 => x"54410083",  4348 => x"78010001",  4349 => x"3c420002",
     4350 => x"38215c90",  4351 => x"b4220800",  4352 => x"28210000",
     4353 => x"c0200000",  4354 => x"29c10000",  4355 => x"b9e01000",
     4356 => x"34030000",  4357 => x"28240014",  4358 => x"15e1001f",
     4359 => x"e0000006",  4360 => x"29c10000",  4361 => x"34020000",
     4362 => x"b9a01800",  4363 => x"28240014",  4364 => x"34010000",
     4365 => x"d8800000",  4366 => x"29610010",  4367 => x"38210002",
     4368 => x"59610010",  4369 => x"e0000057",  4370 => x"296500a8",
     4371 => x"78040001",  4372 => x"b9800800",  4373 => x"34020004",
     4374 => x"34030002",  4375 => x"388442e4",  4376 => x"b9a03000",
     4377 => x"ba003800",  4378 => x"fbfff138",  4379 => x"29c20000",
     4380 => x"296100a8",  4381 => x"28420018",  4382 => x"b6010800",
     4383 => x"596100a8",  4384 => x"d8400000",  4385 => x"29610010",
     4386 => x"38210002",  4387 => x"59610010",  4388 => x"34010005",
     4389 => x"59610014",  4390 => x"e0000058",  4391 => x"78090001",
     4392 => x"39295a38",  4393 => x"29240000",  4394 => x"15e1001f",
     4395 => x"b9e01000",  4396 => x"340300e8",  4397 => x"f80039c1",
     4398 => x"b6027800",  4399 => x"1611001f",  4400 => x"f60f8000",
     4401 => x"b6210800",  4402 => x"b6018000",  4403 => x"15a1001f",
     4404 => x"34030000",  4405 => x"b9a01000",  4406 => x"340403e8",
     4407 => x"f80039b7",  4408 => x"b5e21800",  4409 => x"f5e37800",
     4410 => x"b6010800",  4411 => x"b5e10800",  4412 => x"c8031000",
     4413 => x"48010002",  4414 => x"b8601000",  4415 => x"3401003b",
     4416 => x"4841000d",  4417 => x"29c10000",  4418 => x"34020001",
     4419 => x"28230034",  4420 => x"b9800800",  4421 => x"d8600000",
     4422 => x"296100b0",  4423 => x"59610080",  4424 => x"296100b4",
     4425 => x"59610084",  4426 => x"34010004",  4427 => x"59610014",
     4428 => x"e0000004",  4429 => x"29610088",  4430 => x"34210001",
     4431 => x"59610088",  4432 => x"29620088",  4433 => x"34010009",
     4434 => x"4c22002c",  4435 => x"59600088",  4436 => x"e0000014",
     4437 => x"296300b4",  4438 => x"29610084",  4439 => x"296400b0",
     4440 => x"29620080",  4441 => x"c8610800",  4442 => x"f4231800",
     4443 => x"596100e4",  4444 => x"78010001",  4445 => x"382167c0",
     4446 => x"c8821000",  4447 => x"28210000",  4448 => x"c8431000",
     4449 => x"596200e0",  4450 => x"4420001c",  4451 => x"1601001f",
     4452 => x"34030078",  4453 => x"98301000",  4454 => x"c8411000",
     4455 => x"4c620003",  4456 => x"34010003",  4457 => x"e3ffffbc",
     4458 => x"0021001e",  4459 => x"29c20000",  4460 => x"b4308000",
     4461 => x"296100a8",  4462 => x"16100002",  4463 => x"28420018",
     4464 => x"b6010800",  4465 => x"596100a8",  4466 => x"d8400000",
     4467 => x"296500a8",  4468 => x"78040001",  4469 => x"b9800800",
     4470 => x"34020006",  4471 => x"34030001",  4472 => x"38844300",
     4473 => x"fbfff0d9",  4474 => x"296100b0",  4475 => x"59610080",
     4476 => x"296100b4",  4477 => x"59610084",  4478 => x"29620014",
     4479 => x"34010004",  4480 => x"44410004",  4481 => x"296100f0",
     4482 => x"34210001",  4483 => x"596100f0",  4484 => x"296400e8",
     4485 => x"296300ec",  4486 => x"1481001f",  4487 => x"98611800",
     4488 => x"c8611000",  4489 => x"98812000",  4490 => x"f4431800",
     4491 => x"c8810800",  4492 => x"c8230800",  4493 => x"48200005",
     4494 => x"5c200007",  4495 => x"340101f4",  4496 => x"54410002",
     4497 => x"e0000004",  4498 => x"296100f4",  4499 => x"34210001",
     4500 => x"596100f4",  4501 => x"296500a4",  4502 => x"296400a0",
     4503 => x"ca851800",  4504 => x"f4740800",  4505 => x"cac41000",
     4506 => x"c8411000",  4507 => x"48020007",  4508 => x"34010001",
     4509 => x"48400013",  4510 => x"5c400011",  4511 => x"340203e8",
     4512 => x"54620010",  4513 => x"e000000e",  4514 => x"c8140800",
     4515 => x"7c220000",  4516 => x"c8161800",  4517 => x"c8621800",
     4518 => x"c8251000",  4519 => x"f4410800",  4520 => x"c8641800",
     4521 => x"c8611800",  4522 => x"34010001",  4523 => x"48600005",
     4524 => x"5c600003",  4525 => x"340303e8",  4526 => x"54430002",
     4527 => x"34010000",  4528 => x"202100ff",  4529 => x"44200004",
     4530 => x"296100f8",  4531 => x"34210001",  4532 => x"596100f8",
     4533 => x"78010001",  4534 => x"382192a4",  4535 => x"28210000",
     4536 => x"34020000",  4537 => x"f8000ee2",  4538 => x"29c10000",
     4539 => x"28230038",  4540 => x"44600004",  4541 => x"b9600800",
     4542 => x"34020001",  4543 => x"d8600000",  4544 => x"34010000",
     4545 => x"2b9d0004",  4546 => x"2b8b003c",  4547 => x"2b8c0038",
     4548 => x"2b8d0034",  4549 => x"2b8e0030",  4550 => x"2b8f002c",
     4551 => x"2b900028",  4552 => x"2b910024",  4553 => x"2b920020",
     4554 => x"2b93001c",  4555 => x"2b940018",  4556 => x"2b950014",
     4557 => x"2b960010",  4558 => x"2b97000c",  4559 => x"2b980008",
     4560 => x"379c0044",  4561 => x"c3a00000",  4562 => x"379cffe8",
     4563 => x"5b8b0018",  4564 => x"5b8c0014",  4565 => x"5b8d0010",
     4566 => x"5b8e000c",  4567 => x"5b8f0008",  4568 => x"5b9d0004",
     4569 => x"b8407800",  4570 => x"28220020",  4571 => x"b8205800",
     4572 => x"b8607000",  4573 => x"284d0008",  4574 => x"28220024",
     4575 => x"282c02c8",  4576 => x"28440000",  4577 => x"d8800000",
     4578 => x"48010058",  4579 => x"29610020",  4580 => x"34030008",
     4581 => x"2824000c",  4582 => x"4161004c",  4583 => x"30810004",
     4584 => x"4161004d",  4585 => x"30810005",  4586 => x"4161004e",
     4587 => x"30810006",  4588 => x"3401ffff",  4589 => x"30810007",
     4590 => x"3401fffe",  4591 => x"30810008",  4592 => x"4161004f",
     4593 => x"30810009",  4594 => x"41610050",  4595 => x"3081000a",
     4596 => x"41610051",  4597 => x"3081000b",  4598 => x"29610020",
     4599 => x"2824000c",  4600 => x"b9800800",  4601 => x"34820004",
     4602 => x"f80039c9",  4603 => x"29610020",  4604 => x"35620374",
     4605 => x"28210000",  4606 => x"3180000a",  4607 => x"c8410800",
     4608 => x"14210002",  4609 => x"0821d775",  4610 => x"0d810008",
     4611 => x"41a10042",  4612 => x"3181000b",  4613 => x"34010014",
     4614 => x"3181000c",  4615 => x"41a10043",  4616 => x"3181000d",
     4617 => x"34010002",  4618 => x"3181000e",  4619 => x"78010001",
     4620 => x"3821678c",  4621 => x"28240000",  4622 => x"4480000f",
     4623 => x"b9600800",  4624 => x"b9e01000",  4625 => x"b9c01800",
     4626 => x"d8800000",  4627 => x"4420000a",  4628 => x"78040001",
     4629 => x"78050001",  4630 => x"b9600800",  4631 => x"34020002",
     4632 => x"34030001",  4633 => x"3884436c",  4634 => x"38a55ccc",
     4635 => x"fbfff037",  4636 => x"e000001e",  4637 => x"29610020",
     4638 => x"78040001",  4639 => x"34020003",  4640 => x"2825000c",
     4641 => x"34030001",  4642 => x"b9600800",  4643 => x"40a5000e",
     4644 => x"38844388",  4645 => x"fbfff02d",  4646 => x"29610020",
     4647 => x"78040001",  4648 => x"34020003",  4649 => x"2825000c",
     4650 => x"34030001",  4651 => x"b9600800",  4652 => x"40a5000f",
     4653 => x"3884439c",  4654 => x"fbfff024",  4655 => x"2962003c",
     4656 => x"b9600800",  4657 => x"f8000634",  4658 => x"4162001d",
     4659 => x"34010001",  4660 => x"44410003",  4661 => x"34010004",
     4662 => x"e0000002",  4663 => x"34010006",  4664 => x"59610004",
     4665 => x"e0000003",  4666 => x"340103e8",  4667 => x"59610008",
     4668 => x"34010000",  4669 => x"2b9d0004",  4670 => x"2b8b0018",
     4671 => x"2b8c0014",  4672 => x"2b8d0010",  4673 => x"2b8e000c",
     4674 => x"2b8f0008",  4675 => x"379c0018",  4676 => x"c3a00000",
     4677 => x"379cfff4",  4678 => x"5b8b000c",  4679 => x"5b8c0008",
     4680 => x"5b9d0004",  4681 => x"2822000c",  4682 => x"b8205800",
     4683 => x"44400006",  4684 => x"28220028",  4685 => x"28430018",
     4686 => x"34020fa0",  4687 => x"d8600000",  4688 => x"596102dc",
     4689 => x"296102dc",  4690 => x"44200009",  4691 => x"29610028",
     4692 => x"34020000",  4693 => x"28230018",  4694 => x"b9600800",
     4695 => x"d8600000",  4696 => x"296202dc",  4697 => x"c8220800",
     4698 => x"4c200014",  4699 => x"296c02dc",  4700 => x"34010000",
     4701 => x"4580000a",  4702 => x"29610028",  4703 => x"34020000",
     4704 => x"28230018",  4705 => x"b9600800",  4706 => x"d8600000",
     4707 => x"c9810800",  4708 => x"a4201000",  4709 => x"1442001f",
     4710 => x"a0220800",  4711 => x"59610008",  4712 => x"34010000",
     4713 => x"2b9d0004",  4714 => x"2b8b000c",  4715 => x"2b8c0008",
     4716 => x"379c000c",  4717 => x"c3a00000",  4718 => x"b9600800",
     4719 => x"34020004",  4720 => x"f8000a67",  4721 => x"34010001",
     4722 => x"59610004",  4723 => x"e3fffff5",  4724 => x"340203e8",
     4725 => x"58220008",  4726 => x"34010000",  4727 => x"c3a00000",
     4728 => x"379cfff0",  4729 => x"5b8b0010",  4730 => x"5b8c000c",
     4731 => x"5b8d0008",  4732 => x"5b9d0004",  4733 => x"78040001",
     4734 => x"3884678c",  4735 => x"2884000c",  4736 => x"b8205800",
     4737 => x"b8406800",  4738 => x"b8606000",  4739 => x"44800003",
     4740 => x"d8800000",  4741 => x"5c20001f",  4742 => x"2961000c",
     4743 => x"4420000b",  4744 => x"296102c8",  4745 => x"29630028",
     4746 => x"4022000c",  4747 => x"1021000b",  4748 => x"28630018",
     4749 => x"bc411000",  4750 => x"b9600800",  4751 => x"084203e8",
     4752 => x"d8600000",  4753 => x"596102d4",  4754 => x"4580000f",
     4755 => x"4161030d",  4756 => x"44200008",  4757 => x"3402000b",
     4758 => x"5c22000b",  4759 => x"b9600800",  4760 => x"b9a01000",
     4761 => x"b9801800",  4762 => x"f8000352",  4763 => x"e0000005",
     4764 => x"b9600800",  4765 => x"b9a01000",  4766 => x"b9801800",
     4767 => x"f8000370",  4768 => x"5c200004",  4769 => x"b9600800",
     4770 => x"f800027e",  4771 => x"44200003",  4772 => x"34010002",
     4773 => x"59610004",  4774 => x"29620004",  4775 => x"29610000",
     4776 => x"44410002",  4777 => x"596002d4",  4778 => x"296c02d4",
     4779 => x"34010000",  4780 => x"4580000a",  4781 => x"29610028",
     4782 => x"34020000",  4783 => x"28230018",  4784 => x"b9600800",
     4785 => x"d8600000",  4786 => x"c9810800",  4787 => x"a4201000",
     4788 => x"1442001f",  4789 => x"a0220800",  4790 => x"59610008",
     4791 => x"34010000",  4792 => x"2b9d0004",  4793 => x"2b8b0010",
     4794 => x"2b8c000c",  4795 => x"2b8d0008",  4796 => x"379c0010",
     4797 => x"c3a00000",  4798 => x"34010000",  4799 => x"c3a00000",
     4800 => x"379cffec",  4801 => x"5b8b0014",  4802 => x"5b8c0010",
     4803 => x"5b8d000c",  4804 => x"5b8e0008",  4805 => x"5b9d0004",
     4806 => x"344b00b2",  4807 => x"3d6b0002",  4808 => x"b8407000",
     4809 => x"b42b5800",  4810 => x"29620004",  4811 => x"b8206000",
     4812 => x"340d0000",  4813 => x"44400008",  4814 => x"28220028",
     4815 => x"28430018",  4816 => x"34020000",  4817 => x"d8600000",
     4818 => x"29620004",  4819 => x"c8220800",  4820 => x"4c200009",
     4821 => x"b9a00800",  4822 => x"2b9d0004",  4823 => x"2b8b0014",
     4824 => x"2b8c0010",  4825 => x"2b8d000c",  4826 => x"2b8e0008",
     4827 => x"379c0014",  4828 => x"c3a00000",  4829 => x"b9800800",
     4830 => x"b9c01000",  4831 => x"f80009f8",  4832 => x"340d0001",
     4833 => x"59600004",  4834 => x"e3fffff3",  4835 => x"379cffec",
     4836 => x"5b8b0014",  4837 => x"5b8c0010",  4838 => x"5b8d000c",
     4839 => x"5b8e0008",  4840 => x"5b9d0004",  4841 => x"b8407000",
     4842 => x"2822000c",  4843 => x"b8205800",  4844 => x"b8606800",
     4845 => x"340c0000",  4846 => x"44400014",  4847 => x"282302c8",
     4848 => x"34020001",  4849 => x"1063000d",  4850 => x"f80009f4",
     4851 => x"296302c8",  4852 => x"b9600800",  4853 => x"34020003",
     4854 => x"1063000b",  4855 => x"f80009ef",  4856 => x"29630344",
     4857 => x"34020001",  4858 => x"34010000",  4859 => x"5c620002",
     4860 => x"29610340",  4861 => x"0d61007e",  4862 => x"b9600800",
     4863 => x"f80005d9",  4864 => x"b8206000",  4865 => x"48010047",
     4866 => x"b9600800",  4867 => x"34020001",  4868 => x"fbffffbc",
     4869 => x"44200010",  4870 => x"296302c8",  4871 => x"b9600800",
     4872 => x"34020001",  4873 => x"1063000d",  4874 => x"f80009dc",
     4875 => x"29630344",  4876 => x"34020001",  4877 => x"34010000",
     4878 => x"5c620002",  4879 => x"29610340",  4880 => x"0d61007e",
     4881 => x"b9600800",  4882 => x"f8000613",  4883 => x"48010046",
     4884 => x"340c0000",  4885 => x"b9600800",  4886 => x"34020003",
     4887 => x"fbffffa9",  4888 => x"44200010",  4889 => x"29630344",
     4890 => x"34020001",  4891 => x"34010000",  4892 => x"5c620002",
     4893 => x"29610340",  4894 => x"0d61007e",  4895 => x"b9600800",
     4896 => x"f80005b8",  4897 => x"48010038",  4898 => x"296302c8",
     4899 => x"b9600800",  4900 => x"34020003",  4901 => x"1063000b",
     4902 => x"340c0000",  4903 => x"f80009bf",  4904 => x"45a00020",
     4905 => x"78010001",  4906 => x"3821678c",  4907 => x"28250010",
     4908 => x"4164030d",  4909 => x"44a00007",  4910 => x"b9600800",
     4911 => x"b9c01000",  4912 => x"b9a01800",  4913 => x"d8a00000",
     4914 => x"b8202000",  4915 => x"48010042",  4916 => x"34010001",
     4917 => x"44810010",  4918 => x"3401000b",  4919 => x"44810003",
     4920 => x"5c800010",  4921 => x"e0000006",  4922 => x"b9600800",
     4923 => x"b9c01000",  4924 => x"b9a01800",  4925 => x"f80002af",
     4926 => x"e0000005",  4927 => x"b9600800",  4928 => x"b9c01000",
     4929 => x"b9a01800",  4930 => x"f80002cd",  4931 => x"b8206000",
     4932 => x"e0000004",  4933 => x"b9600800",  4934 => x"356200e4",
     4935 => x"f800066a",  4936 => x"45800006",  4937 => x"34010001",
     4938 => x"4581000f",  4939 => x"3401ffff",  4940 => x"5d81000e",
     4941 => x"e0000029",  4942 => x"29610020",  4943 => x"2821000c",
     4944 => x"4022000e",  4945 => x"340100ff",  4946 => x"44410004",
     4947 => x"4162001d",  4948 => x"34010002",  4949 => x"5c410005",
     4950 => x"34010004",  4951 => x"59610004",  4952 => x"e0000002",
     4953 => x"340c0000",  4954 => x"296e02d8",  4955 => x"340d0000",
     4956 => x"45c0000a",  4957 => x"29610028",  4958 => x"34020000",
     4959 => x"28230018",  4960 => x"b9600800",  4961 => x"d8600000",
     4962 => x"c9c16800",  4963 => x"a5a00800",  4964 => x"1421001f",
     4965 => x"a1a16800",  4966 => x"296e02d0",  4967 => x"34010000",
     4968 => x"45c0000a",  4969 => x"29610028",  4970 => x"34020000",
     4971 => x"28230018",  4972 => x"b9600800",  4973 => x"d8600000",
     4974 => x"c9c10800",  4975 => x"a4201000",  4976 => x"1442001f",
     4977 => x"a0220800",  4978 => x"4da10007",  4979 => x"b9a00800",
     4980 => x"e0000005",  4981 => x"b8206000",  4982 => x"34010002",
     4983 => x"59610004",  4984 => x"340101f4",  4985 => x"59610008",
     4986 => x"b9800800",  4987 => x"2b9d0004",  4988 => x"2b8b0014",
     4989 => x"2b8c0010",  4990 => x"2b8d000c",  4991 => x"2b8e0008",
     4992 => x"379c0014",  4993 => x"c3a00000",  4994 => x"379cfff0",
     4995 => x"5b8b000c",  4996 => x"5b8c0008",  4997 => x"5b9d0004",
     4998 => x"b8406000",  4999 => x"2822000c",  5000 => x"b8205800",
     5001 => x"4440000c",  5002 => x"282202c8",  5003 => x"28250028",
     5004 => x"4044000c",  5005 => x"1042000b",  5006 => x"bc821000",
     5007 => x"28a40018",  5008 => x"084203e8",  5009 => x"5b830010",
     5010 => x"d8800000",  5011 => x"2b830010",  5012 => x"596102d4",
     5013 => x"4460000d",  5014 => x"4161030d",  5015 => x"44200007",
     5016 => x"3402000b",  5017 => x"5c220009",  5018 => x"b9600800",
     5019 => x"b9801000",  5020 => x"f8000250",  5021 => x"e0000004",
     5022 => x"b9600800",  5023 => x"b9801000",  5024 => x"f800026f",
     5025 => x"5c200004",  5026 => x"b9600800",  5027 => x"f800017d",
     5028 => x"44200003",  5029 => x"34010002",  5030 => x"59610004",
     5031 => x"29620004",  5032 => x"29610000",  5033 => x"44410002",
     5034 => x"596002d4",  5035 => x"340103e8",  5036 => x"59610008",
     5037 => x"34010000",  5038 => x"2b9d0004",  5039 => x"2b8b000c",
     5040 => x"2b8c0008",  5041 => x"379c0010",  5042 => x"c3a00000",
     5043 => x"379cfff8",  5044 => x"5b8b0008",  5045 => x"5b9d0004",
     5046 => x"b8205800",  5047 => x"4460000d",  5048 => x"4024030d",
     5049 => x"44800007",  5050 => x"34050008",  5051 => x"44850007",
     5052 => x"3405000b",  5053 => x"5c850007",  5054 => x"f8000198",
     5055 => x"e0000004",  5056 => x"f80001b1",  5057 => x"e0000002",
     5058 => x"f80001e9",  5059 => x"5c200004",  5060 => x"b9600800",
     5061 => x"f800015b",  5062 => x"44200003",  5063 => x"34010002",
     5064 => x"59610004",  5065 => x"340103e8",  5066 => x"59610008",
     5067 => x"34010000",  5068 => x"2b9d0004",  5069 => x"2b8b0008",
     5070 => x"379c0008",  5071 => x"c3a00000",  5072 => x"379cffd4",
     5073 => x"5b8b0014",  5074 => x"5b8c0010",  5075 => x"5b8d000c",
     5076 => x"5b8e0008",  5077 => x"5b9d0004",  5078 => x"b8205800",
     5079 => x"2821000c",  5080 => x"b8407000",  5081 => x"b8606800",
     5082 => x"44200023",  5083 => x"34020000",  5084 => x"34030014",
     5085 => x"35610080",  5086 => x"f8003863",  5087 => x"b9600800",
     5088 => x"f80006da",  5089 => x"78010001",  5090 => x"3821678c",
     5091 => x"28240014",  5092 => x"44800007",  5093 => x"b9600800",
     5094 => x"b9c01000",  5095 => x"b9a01800",  5096 => x"d8800000",
     5097 => x"b8206000",  5098 => x"5c20005f",  5099 => x"4161001c",
     5100 => x"29630028",  5101 => x"202100fd",  5102 => x"3161001c",
     5103 => x"296102c8",  5104 => x"28630018",  5105 => x"4022000c",
     5106 => x"1021000b",  5107 => x"bc411000",  5108 => x"b9600800",
     5109 => x"084203e8",  5110 => x"d8600000",  5111 => x"296302c8",
     5112 => x"596102d4",  5113 => x"34020000",  5114 => x"1063000a",
     5115 => x"b9600800",  5116 => x"f80008ea",  5117 => x"45a00049",
     5118 => x"4161030d",  5119 => x"34020008",  5120 => x"44220012",
     5121 => x"54220003",  5122 => x"5c200044",  5123 => x"e000000a",
     5124 => x"34020009",  5125 => x"44220014",  5126 => x"3402000b",
     5127 => x"5c22003f",  5128 => x"b9600800",  5129 => x"b9c01000",
     5130 => x"b9a01800",  5131 => x"f800014b",  5132 => x"e000000a",
     5133 => x"b9600800",  5134 => x"b9c01000",  5135 => x"b9a01800",
     5136 => x"f8000161",  5137 => x"e0000005",  5138 => x"b9600800",
     5139 => x"b9c01000",  5140 => x"b9a01800",  5141 => x"f8000196",
     5142 => x"b8206000",  5143 => x"5c200032",  5144 => x"e000002e",
     5145 => x"34010035",  5146 => x"340c0001",  5147 => x"4c2d002e",
     5148 => x"378c0018",  5149 => x"b9c00800",  5150 => x"b9801000",
     5151 => x"f80004a2",  5152 => x"296102c8",  5153 => x"37820024",
     5154 => x"34030008",  5155 => x"f800377f",  5156 => x"5c20001c",
     5157 => x"2d6202f2",  5158 => x"2d61032a",  5159 => x"5c410019",
     5160 => x"296102c8",  5161 => x"2c220008",  5162 => x"2f81002c",
     5163 => x"5c410015",  5164 => x"4161001c",  5165 => x"20210001",
     5166 => x"44200012",  5167 => x"b9801000",  5168 => x"356100bc",
     5169 => x"f8000619",  5170 => x"78010001",  5171 => x"3821678c",
     5172 => x"28220018",  5173 => x"44400006",  5174 => x"b9600800",
     5175 => x"d8400000",  5176 => x"b8206000",  5177 => x"5c200010",
     5178 => x"e0000003",  5179 => x"b9600800",  5180 => x"f80006d7",
     5181 => x"4161032d",  5182 => x"316102ee",  5183 => x"e0000007",
     5184 => x"78040001",  5185 => x"b9600800",  5186 => x"34020005",
     5187 => x"34030002",  5188 => x"388443b4",  5189 => x"fbffee0d",
     5190 => x"b9600800",  5191 => x"f80000d9",  5192 => x"b8206000",
     5193 => x"296102cc",  5194 => x"44200009",  5195 => x"29610028",
     5196 => x"34020000",  5197 => x"28230018",  5198 => x"b9600800",
     5199 => x"d8600000",  5200 => x"296202cc",  5201 => x"c8220800",
     5202 => x"4c200033",  5203 => x"3401ffff",  5204 => x"45810005",
     5205 => x"7d810001",  5206 => x"c8010800",  5207 => x"a1816000",
     5208 => x"e0000003",  5209 => x"34010002",  5210 => x"59610004",
     5211 => x"29620004",  5212 => x"29610000",  5213 => x"44410005",
     5214 => x"596002d4",  5215 => x"596002cc",  5216 => x"b9600800",
     5217 => x"f8000659",  5218 => x"296e02d4",  5219 => x"340d0000",
     5220 => x"45c0000a",  5221 => x"29610028",  5222 => x"34020000",
     5223 => x"28230018",  5224 => x"b9600800",  5225 => x"d8600000",
     5226 => x"c9c16800",  5227 => x"a5a00800",  5228 => x"1421001f",
     5229 => x"a1a16800",  5230 => x"296e02cc",  5231 => x"b9a00800",
     5232 => x"45c0000a",  5233 => x"29610028",  5234 => x"34020000",
     5235 => x"28230018",  5236 => x"b9600800",  5237 => x"d8600000",
     5238 => x"c9c10800",  5239 => x"a4201000",  5240 => x"1442001f",
     5241 => x"a0220800",  5242 => x"4da10002",  5243 => x"b9a00800",
     5244 => x"59610008",  5245 => x"b9800800",  5246 => x"2b9d0004",
     5247 => x"2b8b0014",  5248 => x"2b8c0010",  5249 => x"2b8d000c",
     5250 => x"2b8e0008",  5251 => x"379c002c",  5252 => x"c3a00000",
     5253 => x"b9600800",  5254 => x"34020000",  5255 => x"f8000850",
     5256 => x"b9600800",  5257 => x"596002cc",  5258 => x"f80004f6",
     5259 => x"29630100",  5260 => x"29620104",  5261 => x"296500f8",
     5262 => x"296400fc",  5263 => x"b8206000",  5264 => x"29610108",
     5265 => x"596300b0",  5266 => x"296302c8",  5267 => x"596200b4",
     5268 => x"596100b8",  5269 => x"596500a8",  5270 => x"596400ac",
     5271 => x"1063000a",  5272 => x"b9600800",  5273 => x"34020000",
     5274 => x"f800084c",  5275 => x"29620020",  5276 => x"356100a8",
     5277 => x"28430008",  5278 => x"b8201000",  5279 => x"34630018",
     5280 => x"f80005bd",  5281 => x"e3ffffb2",  5282 => x"379cfff8",
     5283 => x"5b8b0008",  5284 => x"5b9d0004",  5285 => x"282202c8",
     5286 => x"28240028",  5287 => x"b8205800",  5288 => x"4043000c",
     5289 => x"1042000b",  5290 => x"bc621000",  5291 => x"28830018",
     5292 => x"084203e8",  5293 => x"d8600000",  5294 => x"596102d4",
     5295 => x"2b9d0004",  5296 => x"2b8b0008",  5297 => x"379c0008",
     5298 => x"c3a00000",  5299 => x"379cffe4",  5300 => x"5b8b001c",
     5301 => x"5b8c0018",  5302 => x"5b8d0014",  5303 => x"5b8e0010",
     5304 => x"5b8f000c",  5305 => x"5b900008",  5306 => x"5b9d0004",
     5307 => x"340c0000",  5308 => x"b8205800",  5309 => x"b8407000",
     5310 => x"342f030c",  5311 => x"34300320",  5312 => x"e0000013",
     5313 => x"098d0058",  5314 => x"ba000800",  5315 => x"3403000a",
     5316 => x"35a20110",  5317 => x"b5621000",  5318 => x"f80036dc",
     5319 => x"5c20000b",  5320 => x"b56d0800",  5321 => x"b9e01000",
     5322 => x"34030024",  5323 => x"34210144",  5324 => x"f80036f7",
     5325 => x"b56d5800",  5326 => x"b9c00800",  5327 => x"3562011c",
     5328 => x"f80003be",  5329 => x"e0000020",  5330 => x"358c0001",
     5331 => x"2d63010c",  5332 => x"486cffed",  5333 => x"34010004",
     5334 => x"54610003",  5335 => x"34630001",  5336 => x"0d63010c",
     5337 => x"2d6d010c",  5338 => x"35620320",  5339 => x"3403000a",
     5340 => x"35adffff",  5341 => x"09ac0058",  5342 => x"35810110",
     5343 => x"b5610800",  5344 => x"f80036e3",  5345 => x"b56c0800",
     5346 => x"34030024",  5347 => x"b9e01000",  5348 => x"34210144",
     5349 => x"f80036de",  5350 => x"b56c1000",  5351 => x"b9c00800",
     5352 => x"3442011c",  5353 => x"f80003a5",  5354 => x"78040001",
     5355 => x"b9600800",  5356 => x"34020003",  5357 => x"34030001",
     5358 => x"388443e4",  5359 => x"b9a02800",  5360 => x"fbffed62",
     5361 => x"2b9d0004",  5362 => x"2b8b001c",  5363 => x"2b8c0018",
     5364 => x"2b8d0014",  5365 => x"2b8e0010",  5366 => x"2b8f000c",
     5367 => x"2b900008",  5368 => x"379c001c",  5369 => x"c3a00000",
     5370 => x"4022001e",  5371 => x"34030001",  5372 => x"44430009",
     5373 => x"44400008",  5374 => x"34030002",  5375 => x"5c430008",
     5376 => x"34020012",  5377 => x"58220070",  5378 => x"3402000e",
     5379 => x"58220074",  5380 => x"e0000003",  5381 => x"58200070",
     5382 => x"58200074",  5383 => x"28240070",  5384 => x"2825002c",
     5385 => x"34020000",  5386 => x"b4a42800",  5387 => x"20a30003",
     5388 => x"44600003",  5389 => x"34020004",  5390 => x"c8431000",
     5391 => x"b4a22800",  5392 => x"28260030",  5393 => x"28220074",
     5394 => x"5825003c",  5395 => x"34030000",  5396 => x"b4c23000",
     5397 => x"20c70003",  5398 => x"44e00003",  5399 => x"34030004",
     5400 => x"c8671800",  5401 => x"b4c31800",  5402 => x"c8a42000",
     5403 => x"c8621000",  5404 => x"58230040",  5405 => x"58240034",
     5406 => x"58220038",  5407 => x"c3a00000",  5408 => x"379cfff4",
     5409 => x"5b8b000c",  5410 => x"5b8c0008",  5411 => x"5b9d0004",
     5412 => x"78020001",  5413 => x"3842678c",  5414 => x"28420020",
     5415 => x"b8205800",  5416 => x"44400006",  5417 => x"d8400000",
     5418 => x"b8206000",  5419 => x"34010001",  5420 => x"45810018",
     5421 => x"480c0018",  5422 => x"296102d4",  5423 => x"340c0000",
     5424 => x"44200015",  5425 => x"29610028",  5426 => x"34020000",
     5427 => x"28230018",  5428 => x"b9600800",  5429 => x"d8600000",
     5430 => x"296202d4",  5431 => x"c8220800",  5432 => x"4c200013",
     5433 => x"e000000c",  5434 => x"4162001d",  5435 => x"34010002",
     5436 => x"44410004",  5437 => x"34010006",  5438 => x"59610004",
     5439 => x"e0000006",  5440 => x"34010004",  5441 => x"59610004",
     5442 => x"b9600800",  5443 => x"fbffff5f",  5444 => x"340c0000",
     5445 => x"b9800800",  5446 => x"2b9d0004",  5447 => x"2b8b000c",
     5448 => x"2b8c0008",  5449 => x"379c000c",  5450 => x"c3a00000",
     5451 => x"b9600800",  5452 => x"34020002",  5453 => x"f800078a",
     5454 => x"29610020",  5455 => x"596002d4",  5456 => x"0d60010c",
     5457 => x"2821000c",  5458 => x"4022000e",  5459 => x"340100ff",
     5460 => x"5c41ffe6",  5461 => x"e3ffffeb",  5462 => x"379cfff4",
     5463 => x"5b8b000c",  5464 => x"5b8c0008",  5465 => x"5b9d0004",
     5466 => x"3404003f",  5467 => x"b8205800",  5468 => x"340cffff",
     5469 => x"4c83000e",  5470 => x"fbffff55",  5471 => x"b9600800",
     5472 => x"fbffff42",  5473 => x"b9600800",  5474 => x"f800015a",
     5475 => x"59610004",  5476 => x"78010001",  5477 => x"3821678c",
     5478 => x"28220024",  5479 => x"340c0000",  5480 => x"44400003",
     5481 => x"b9600800",  5482 => x"d8400000",  5483 => x"b9800800",
     5484 => x"2b9d0004",  5485 => x"2b8b000c",  5486 => x"2b8c0008",
     5487 => x"379c000c",  5488 => x"c3a00000",  5489 => x"379cffe0",
     5490 => x"5b8b0014",  5491 => x"5b8c0010",  5492 => x"5b8d000c",
     5493 => x"5b8e0008",  5494 => x"5b9d0004",  5495 => x"b8205800",
     5496 => x"3401002b",  5497 => x"b8407000",  5498 => x"340cffff",
     5499 => x"4c230028",  5500 => x"4161001c",  5501 => x"340c0000",
     5502 => x"20210001",  5503 => x"44200024",  5504 => x"296300ec",
     5505 => x"296200f0",  5506 => x"296100f4",  5507 => x"296500e4",
     5508 => x"296400e8",  5509 => x"5963009c",  5510 => x"596200a0",
     5511 => x"2963031c",  5512 => x"29620318",  5513 => x"596100a4",
     5514 => x"59650094",  5515 => x"356100d0",  5516 => x"59640098",
     5517 => x"f8000485",  5518 => x"41610313",  5519 => x"20210002",
     5520 => x"44200007",  5521 => x"4161001c",  5522 => x"38210002",
     5523 => x"3161001c",  5524 => x"2d61032a",  5525 => x"0d6102ec",
     5526 => x"e000000d",  5527 => x"378d0018",  5528 => x"b9c00800",
     5529 => x"b9a01000",  5530 => x"f80002ed",  5531 => x"4161001c",
     5532 => x"b9a01000",  5533 => x"202100fd",  5534 => x"3161001c",
     5535 => x"35610080",  5536 => x"f80004aa",  5537 => x"b9600800",
     5538 => x"f8000551",  5539 => x"b9800800",  5540 => x"2b9d0004",
     5541 => x"2b8b0014",  5542 => x"2b8c0010",  5543 => x"2b8d000c",
     5544 => x"2b8e0008",  5545 => x"379c0020",  5546 => x"c3a00000",
     5547 => x"379cffe4",  5548 => x"5b8b0010",  5549 => x"5b8c000c",
     5550 => x"5b8d0008",  5551 => x"5b9d0004",  5552 => x"b8205800",
     5553 => x"b8400800",  5554 => x"3402002b",  5555 => x"3404ffff",
     5556 => x"4c430031",  5557 => x"4162001c",  5558 => x"20430001",
     5559 => x"5c600004",  5560 => x"78010001",  5561 => x"38214404",
     5562 => x"e0000005",  5563 => x"20420002",  5564 => x"5c400007",
     5565 => x"78010001",  5566 => x"38214440",  5567 => x"78020001",
     5568 => x"38425cdc",  5569 => x"f8001c2e",  5570 => x"e0000022",
     5571 => x"2d6402ec",  5572 => x"2d63032a",  5573 => x"44830007",
     5574 => x"78010001",  5575 => x"78020001",  5576 => x"38425cdc",
     5577 => x"38214478",  5578 => x"f8001c25",  5579 => x"e0000019",
     5580 => x"378d0014",  5581 => x"b9a01000",  5582 => x"f80002ec",
     5583 => x"4161001c",  5584 => x"356c0080",  5585 => x"b9a01000",
     5586 => x"202100fd",  5587 => x"3161001c",  5588 => x"b9800800",
     5589 => x"f8000475",  5590 => x"78030001",  5591 => x"3863678c",
     5592 => x"28640028",  5593 => x"44800009",  5594 => x"b9600800",
     5595 => x"b9801000",  5596 => x"356300d0",  5597 => x"d8800000",
     5598 => x"b8202000",  5599 => x"34010001",  5600 => x"44810004",
     5601 => x"48040004",  5602 => x"b9600800",  5603 => x"f8000510",
     5604 => x"34040000",  5605 => x"b8800800",  5606 => x"2b9d0004",
     5607 => x"2b8b0010",  5608 => x"2b8c000c",  5609 => x"2b8d0008",
     5610 => x"379c001c",  5611 => x"c3a00000",  5612 => x"379cfff0",
     5613 => x"5b8b0010",  5614 => x"5b8c000c",  5615 => x"5b8d0008",
     5616 => x"5b9d0004",  5617 => x"b8406800",  5618 => x"3402003f",
     5619 => x"b8205800",  5620 => x"340cffff",  5621 => x"4c430013",
     5622 => x"78040001",  5623 => x"34030002",  5624 => x"388444b8",
     5625 => x"34020003",  5626 => x"fbffec58",  5627 => x"b9a01000",
     5628 => x"b9600800",  5629 => x"fbfffeb6",  5630 => x"b9600800",
     5631 => x"f80000bd",  5632 => x"59610004",  5633 => x"78010001",
     5634 => x"3821678c",  5635 => x"28220024",  5636 => x"340c0000",
     5637 => x"44400003",  5638 => x"b9600800",  5639 => x"d8400000",
     5640 => x"b9800800",  5641 => x"2b9d0004",  5642 => x"2b8b0010",
     5643 => x"2b8c000c",  5644 => x"2b8d0008",  5645 => x"379c0010",
     5646 => x"c3a00000",  5647 => x"34010000",  5648 => x"c3a00000",
     5649 => x"379cfffc",  5650 => x"5b9d0004",  5651 => x"34030008",
     5652 => x"f800358e",  5653 => x"2b9d0004",  5654 => x"379c0004",
     5655 => x"c3a00000",  5656 => x"379cffe0",  5657 => x"5b8b0020",
     5658 => x"5b8c001c",  5659 => x"5b8d0018",  5660 => x"5b8e0014",
     5661 => x"5b8f0010",  5662 => x"5b90000c",  5663 => x"5b910008",
     5664 => x"5b9d0004",  5665 => x"780e0001",  5666 => x"39ce5cfc",
     5667 => x"78040001",  5668 => x"b8406800",  5669 => x"b8606000",
     5670 => x"34020003",  5671 => x"34030002",  5672 => x"38844860",
     5673 => x"b9c02800",  5674 => x"b8207800",  5675 => x"35b10021",
     5676 => x"fbffec26",  5677 => x"35900021",  5678 => x"ba200800",
     5679 => x"ba001000",  5680 => x"fbffffe1",  5681 => x"5c200033",
     5682 => x"2d81002a",  5683 => x"2dab002a",  5684 => x"c9615800",
     5685 => x"35620001",  5686 => x"34010002",  5687 => x"54410043",
     5688 => x"29e20020",  5689 => x"34030001",  5690 => x"35a10048",
     5691 => x"28420014",  5692 => x"5d63000b",  5693 => x"fbffffd4",
     5694 => x"5c20003c",  5695 => x"78040001",  5696 => x"b9e00800",
     5697 => x"34020003",  5698 => x"34030001",  5699 => x"388444e8",
     5700 => x"b9c02800",  5701 => x"3406008f",  5702 => x"e000000e",
     5703 => x"3403ffff",  5704 => x"358c0048",  5705 => x"5d63000e",
     5706 => x"b9800800",  5707 => x"fbffffc6",  5708 => x"5c20002e",
     5709 => x"78040001",  5710 => x"b9e00800",  5711 => x"34020003",
     5712 => x"34030001",  5713 => x"388444e8",  5714 => x"b9c02800",
     5715 => x"34060098",  5716 => x"fbffebfe",  5717 => x"340b0000",
     5718 => x"e0000024",  5719 => x"b9801000",  5720 => x"fbffffb9",
     5721 => x"b8205800",  5722 => x"5c200020",  5723 => x"78040001",
     5724 => x"b9e00800",  5725 => x"34020003",  5726 => x"34030001",
     5727 => x"388444f8",  5728 => x"b9c02800",  5729 => x"340600a0",
     5730 => x"fbffebf0",  5731 => x"e0000017",  5732 => x"41ab001a",
     5733 => x"4181001a",  5734 => x"5d61000e",  5735 => x"41ab001c",
     5736 => x"4181001c",  5737 => x"5d61000b",  5738 => x"41ab001d",
     5739 => x"4181001d",  5740 => x"5d610008",  5741 => x"2da2001e",
     5742 => x"2d81001e",  5743 => x"340b0000",  5744 => x"5c41000a",
     5745 => x"41ab0020",  5746 => x"41810020",  5747 => x"45610003",
     5748 => x"c9615800",  5749 => x"e0000005",  5750 => x"ba200800",
     5751 => x"ba001000",  5752 => x"fbffff99",  5753 => x"b8205800",
     5754 => x"b9600800",  5755 => x"2b9d0004",  5756 => x"2b8b0020",
     5757 => x"2b8c001c",  5758 => x"2b8d0018",  5759 => x"2b8e0014",
     5760 => x"2b8f0010",  5761 => x"2b90000c",  5762 => x"2b910008",
     5763 => x"379c0020",  5764 => x"c3a00000",  5765 => x"379cfffc",
     5766 => x"5b9d0004",  5767 => x"34020000",  5768 => x"34030014",
     5769 => x"f80035b8",  5770 => x"2b9d0004",  5771 => x"379c0004",
     5772 => x"c3a00000",  5773 => x"379cfff0",  5774 => x"5b8b0010",
     5775 => x"5b8c000c",  5776 => x"5b8d0008",  5777 => x"5b9d0004",
     5778 => x"b8206800",  5779 => x"28210020",  5780 => x"282c0014",
     5781 => x"282b000c",  5782 => x"28210010",  5783 => x"0c200000",
     5784 => x"34210004",  5785 => x"fbffffec",  5786 => x"29a10020",
     5787 => x"28210010",  5788 => x"34210018",  5789 => x"fbffffe8",
     5790 => x"b9800800",  5791 => x"34020000",  5792 => x"34030020",
     5793 => x"f80035a0",  5794 => x"29610004",  5795 => x"3402ffa0",
     5796 => x"59810000",  5797 => x"29610008",  5798 => x"59810004",
     5799 => x"29610004",  5800 => x"59810010",  5801 => x"29610008",
     5802 => x"59810014",  5803 => x"2d61000e",  5804 => x"0d810018",
     5805 => x"2d610010",  5806 => x"0d81001a",  5807 => x"41610012",
     5808 => x"3181001c",  5809 => x"41610013",  5810 => x"3181001d",
     5811 => x"29a10020",  5812 => x"28210018",  5813 => x"3022001c",
     5814 => x"2b9d0004",  5815 => x"2b8b0010",  5816 => x"2b8c000c",
     5817 => x"2b8d0008",  5818 => x"379c0010",  5819 => x"c3a00000",
     5820 => x"379cff8c",  5821 => x"5b8b0018",  5822 => x"5b8c0014",
     5823 => x"5b8d0010",  5824 => x"5b8e000c",  5825 => x"5b8f0008",
     5826 => x"5b9d0004",  5827 => x"2c22010c",  5828 => x"b8205800",
     5829 => x"340d0000",  5830 => x"340c0001",  5831 => x"5c400014",
     5832 => x"28230000",  5833 => x"b8406800",  5834 => x"34020006",
     5835 => x"5c620010",  5836 => x"fbffffc1",  5837 => x"29610000",
     5838 => x"e0000105",  5839 => x"09820058",  5840 => x"09a30058",
     5841 => x"b9600800",  5842 => x"34420110",  5843 => x"34630110",
     5844 => x"b5621000",  5845 => x"b5631800",  5846 => x"fbffff42",
     5847 => x"48010002",  5848 => x"e0000002",  5849 => x"b9806800",
     5850 => x"358c0001",  5851 => x"2d66010c",  5852 => x"48ccfff3",
     5853 => x"78040001",  5854 => x"b9600800",  5855 => x"34020003",
     5856 => x"34030001",  5857 => x"38844508",  5858 => x"b9a02800",
     5859 => x"fbffeb6f",  5860 => x"1d61010e",  5861 => x"442d0022",
     5862 => x"0d6d010e",  5863 => x"296c0020",  5864 => x"340f0000",
     5865 => x"340e0001",  5866 => x"e0000015",  5867 => x"29820000",
     5868 => x"09c10374",  5869 => x"b4410800",  5870 => x"2c23010c",
     5871 => x"4460000f",  5872 => x"09e40374",  5873 => x"1c23010e",
     5874 => x"b4442000",  5875 => x"1c82010e",  5876 => x"08630058",
     5877 => x"08420058",  5878 => x"34630110",  5879 => x"b4231800",
     5880 => x"34420110",  5881 => x"b4821000",  5882 => x"fbffff1e",
     5883 => x"48010002",  5884 => x"e0000002",  5885 => x"b9c07800",
     5886 => x"35ce0001",  5887 => x"2981000c",  5888 => x"2c21000c",
     5889 => x"482effea",  5890 => x"2981001c",  5891 => x"442f0004",
     5892 => x"34010001",  5893 => x"598f001c",  5894 => x"59810020",
     5895 => x"4162001d",  5896 => x"34010002",  5897 => x"44410063",
     5898 => x"2d61010c",  5899 => x"5c200004",  5900 => x"29620000",
     5901 => x"34010004",  5902 => x"444100c5",  5903 => x"29610020",
     5904 => x"09ac0058",  5905 => x"2821000c",  5906 => x"4023000a",
     5907 => x"4022000b",  5908 => x"40290004",  5909 => x"40280005",
     5910 => x"40270006",  5911 => x"40260007",  5912 => x"40250008",
     5913 => x"40240009",  5914 => x"33830047",  5915 => x"33890041",
     5916 => x"33880042",  5917 => x"33870043",  5918 => x"33860044",
     5919 => x"33850045",  5920 => x"33840046",  5921 => x"33820048",
     5922 => x"2c22000e",  5923 => x"35830110",  5924 => x"b5631800",
     5925 => x"0f82003c",  5926 => x"2c220010",  5927 => x"0f82003e",
     5928 => x"40220012",  5929 => x"3382003a",  5930 => x"40220013",
     5931 => x"0f80004a",  5932 => x"33820040",  5933 => x"28220004",
     5934 => x"5b820068",  5935 => x"28210008",  5936 => x"37820020",
     5937 => x"5b81006c",  5938 => x"b9600800",  5939 => x"fbfffee5",
     5940 => x"4162001d",  5941 => x"34030001",  5942 => x"44430029",
     5943 => x"29620020",  5944 => x"78050001",  5945 => x"38a55d0c",
     5946 => x"2844000c",  5947 => x"1086000e",  5948 => x"48060004",
     5949 => x"48010023",  5950 => x"5c200019",  5951 => x"e0000006",
     5952 => x"48010020",  5953 => x"44200004",  5954 => x"2c81000c",
     5955 => x"5c23000a",  5956 => x"e0000028",  5957 => x"78040001",
     5958 => x"b9600800",  5959 => x"34020003",  5960 => x"34030001",
     5961 => x"38844528",  5962 => x"fbffeb08",  5963 => x"34010002",
     5964 => x"e0000087",  5965 => x"29630338",  5966 => x"2841001c",
     5967 => x"4461001d",  5968 => x"b56c1000",  5969 => x"37810041",
     5970 => x"34420131",  5971 => x"5b85001c",  5972 => x"fbfffebd",
     5973 => x"2b85001c",  5974 => x"5c20000c",  5975 => x"78040001",
     5976 => x"b9600800",  5977 => x"34020003",  5978 => x"34030001",
     5979 => x"38844534",  5980 => x"fbffeaf6",  5981 => x"34010007",
     5982 => x"e0000075",  5983 => x"4c200003",  5984 => x"b9600800",
     5985 => x"fbffff2c",  5986 => x"78040001",  5987 => x"78050001",
     5988 => x"b9600800",  5989 => x"34020003",  5990 => x"34030001",
     5991 => x"38844544",  5992 => x"38a55d0c",  5993 => x"fbffeae9",
     5994 => x"34010006",  5995 => x"e0000068",  5996 => x"09a30058",
     5997 => x"29620020",  5998 => x"b5631800",  5999 => x"2c64013a",
     6000 => x"284c0018",  6001 => x"28410014",  6002 => x"28420010",
     6003 => x"34840001",  6004 => x"0c440000",  6005 => x"34620150",
     6006 => x"28450008",  6007 => x"2844000c",  6008 => x"58250000",
     6009 => x"58240004",  6010 => x"2c420010",  6011 => x"0c220008",
     6012 => x"34620128",  6013 => x"404e0009",  6014 => x"4045000f",
     6015 => x"40440010",  6016 => x"404a000a",  6017 => x"4049000b",
     6018 => x"4048000c",  6019 => x"4047000d",  6020 => x"4046000e",
     6021 => x"302e0010",  6022 => x"30250016",  6023 => x"302a0011",
     6024 => x"30290012",  6025 => x"30280013",  6026 => x"30270014",
     6027 => x"30260015",  6028 => x"30240017",  6029 => x"28440004",
     6030 => x"346e0120",  6031 => x"58240018",  6032 => x"41c4000a",
     6033 => x"3024001c",  6034 => x"40420008",  6035 => x"3022001d",
     6036 => x"4061013c",  6037 => x"3181001c",  6038 => x"1dc50008",
     6039 => x"1d810000",  6040 => x"4425000e",  6041 => x"78040001",
     6042 => x"b9600800",  6043 => x"34020003",  6044 => x"34030001",
     6045 => x"38844550",  6046 => x"fbffeab4",  6047 => x"2dc10008",
     6048 => x"34020000",  6049 => x"0d810000",  6050 => x"29610028",
     6051 => x"28230004",  6052 => x"b9600800",  6053 => x"d8600000",
     6054 => x"09ad0058",  6055 => x"b56d0800",  6056 => x"34210141",
     6057 => x"4022000b",  6058 => x"20420004",  6059 => x"7c420000",
     6060 => x"59820004",  6061 => x"4022000b",  6062 => x"20420002",
     6063 => x"7c420000",  6064 => x"59820008",  6065 => x"4022000b",
     6066 => x"20420001",  6067 => x"5982000c",  6068 => x"4022000b",
     6069 => x"20420010",  6070 => x"7c420000",  6071 => x"59820010",
     6072 => x"4022000b",  6073 => x"20420020",  6074 => x"7c420000",
     6075 => x"59820014",  6076 => x"4021000b",  6077 => x"20210008",
     6078 => x"7c210000",  6079 => x"59810018",  6080 => x"78010001",
     6081 => x"3821678c",  6082 => x"2824001c",  6083 => x"44800007",
     6084 => x"b56d1000",  6085 => x"b8406800",  6086 => x"b9600800",
     6087 => x"34420144",  6088 => x"35a3011c",  6089 => x"d8800000",
     6090 => x"78040001",  6091 => x"78050001",  6092 => x"b9600800",
     6093 => x"34020003",  6094 => x"34030001",  6095 => x"38844564",
     6096 => x"38a55d0c",  6097 => x"fbffea81",  6098 => x"34010009",
     6099 => x"2b9d0004",  6100 => x"2b8b0018",  6101 => x"2b8c0014",
     6102 => x"2b8d0010",  6103 => x"2b8e000c",  6104 => x"2b8f0008",
     6105 => x"379c0074",  6106 => x"c3a00000",  6107 => x"379cffec",
     6108 => x"5b8b0014",  6109 => x"5b8c0010",  6110 => x"5b8d000c",
     6111 => x"5b8e0008",  6112 => x"5b9d0004",  6113 => x"b8406000",
     6114 => x"28220024",  6115 => x"b8607000",  6116 => x"28230070",
     6117 => x"2847000c",  6118 => x"28220034",  6119 => x"b8806800",
     6120 => x"b5831800",  6121 => x"342400f8",  6122 => x"b9a02800",
     6123 => x"34060000",  6124 => x"b8205800",  6125 => x"d8e00000",
     6126 => x"78070001",  6127 => x"38e767c4",  6128 => x"3dc20002",
     6129 => x"4c2c000c",  6130 => x"b4e23800",  6131 => x"28e50000",
     6132 => x"78040001",  6133 => x"b9600800",  6134 => x"34020005",
     6135 => x"34030001",  6136 => x"3884419c",  6137 => x"b9c03000",
     6138 => x"fbffea58",  6139 => x"3401ffff",  6140 => x"e0000014",
     6141 => x"b4e24000",  6142 => x"296600f8",  6143 => x"296700fc",
     6144 => x"29080000",  6145 => x"78040001",  6146 => x"b9600800",
     6147 => x"34020005",  6148 => x"34030001",  6149 => x"388441bc",
     6150 => x"b9802800",  6151 => x"fbffea4b",  6152 => x"34010001",
     6153 => x"5da10003",  6154 => x"29620104",  6155 => x"44400005",
     6156 => x"2961036c",  6157 => x"34210001",  6158 => x"5961036c",
     6159 => x"34010000",  6160 => x"2b9d0004",  6161 => x"2b8b0014",
     6162 => x"2b8c0010",  6163 => x"2b8d000c",  6164 => x"2b8e0008",
     6165 => x"379c0014",  6166 => x"c3a00000",  6167 => x"379cfff0",
     6168 => x"5b8b0010",  6169 => x"5b8c000c",  6170 => x"5b8d0008",
     6171 => x"5b9d0004",  6172 => x"b8205800",  6173 => x"40410000",
     6174 => x"b8406000",  6175 => x"34030002",  6176 => x"00210004",
     6177 => x"356d0320",  6178 => x"3161030c",  6179 => x"40410000",
     6180 => x"2021000f",  6181 => x"3161030d",  6182 => x"40410001",
     6183 => x"2021000f",  6184 => x"3161030e",  6185 => x"2c410002",
     6186 => x"0d610310",  6187 => x"40410004",  6188 => x"34420006",
     6189 => x"31610312",  6190 => x"35610313",  6191 => x"f8003394",
     6192 => x"35820008",  6193 => x"34030004",  6194 => x"3561031c",
     6195 => x"f8003390",  6196 => x"3582000c",  6197 => x"34030004",
     6198 => x"35610318",  6199 => x"f800338c",  6200 => x"35820014",
     6201 => x"34030008",  6202 => x"b9a00800",  6203 => x"f8003388",
     6204 => x"2d81001c",  6205 => x"296202c8",  6206 => x"34030008",
     6207 => x"0d610328",  6208 => x"2d81001e",  6209 => x"0d61032a",
     6210 => x"41810020",  6211 => x"3161032c",  6212 => x"41810021",
     6213 => x"3161032d",  6214 => x"b9a00800",  6215 => x"f800335b",
     6216 => x"3403ffff",  6217 => x"44200015",  6218 => x"29610020",
     6219 => x"28210014",  6220 => x"2c220008",  6221 => x"4440000a",
     6222 => x"b9a01000",  6223 => x"34030008",  6224 => x"f8003352",
     6225 => x"5c200009",  6226 => x"29610020",  6227 => x"28210014",
     6228 => x"2c220008",  6229 => x"2d610328",  6230 => x"5c410004",
     6231 => x"4161001c",  6232 => x"38210001",  6233 => x"e0000003",
     6234 => x"4161001c",  6235 => x"202100fe",  6236 => x"3161001c",
     6237 => x"34030000",  6238 => x"b8600800",  6239 => x"2b9d0004",
     6240 => x"2b8b0010",  6241 => x"2b8c000c",  6242 => x"2b8d0008",
     6243 => x"379c0010",  6244 => x"c3a00000",  6245 => x"379cfff4",
     6246 => x"5b8b000c",  6247 => x"5b8c0008",  6248 => x"5b9d0004",
     6249 => x"30400000",  6250 => x"b8206000",  6251 => x"282102c8",
     6252 => x"b8405800",  6253 => x"34030008",  6254 => x"4021000e",
     6255 => x"30410001",  6256 => x"29810020",  6257 => x"2821000c",
     6258 => x"40210014",  6259 => x"30410004",  6260 => x"34010002",
     6261 => x"30410006",  6262 => x"34410008",  6263 => x"34020000",
     6264 => x"f80033c9",  6265 => x"298202c8",  6266 => x"35610014",
     6267 => x"34030008",  6268 => x"f8003347",  6269 => x"298102c8",
     6270 => x"2c210008",  6271 => x"0d61001c",  6272 => x"3401007f",
     6273 => x"31610021",  6274 => x"2b9d0004",  6275 => x"2b8b000c",
     6276 => x"2b8c0008",  6277 => x"379c000c",  6278 => x"c3a00000",
     6279 => x"2c230022",  6280 => x"0c430004",  6281 => x"28230024",
     6282 => x"58430000",  6283 => x"28210028",  6284 => x"58410008",
     6285 => x"c3a00000",  6286 => x"379cfff4",  6287 => x"5b8b000c",
     6288 => x"5b8c0008",  6289 => x"5b9d0004",  6290 => x"b8205800",
     6291 => x"2c210022",  6292 => x"b8406000",  6293 => x"34030008",
     6294 => x"0c410004",  6295 => x"29610024",  6296 => x"58410000",
     6297 => x"29610028",  6298 => x"58410008",  6299 => x"2d61002c",
     6300 => x"0c41000c",  6301 => x"4161002f",  6302 => x"3041000e",
     6303 => x"41610030",  6304 => x"30410010",  6305 => x"41610031",
     6306 => x"30410011",  6307 => x"2d610032",  6308 => x"0c410012",
     6309 => x"41610034",  6310 => x"30410014",  6311 => x"34410015",
     6312 => x"35620035",  6313 => x"f800331a",  6314 => x"2d61003d",
     6315 => x"0d81001e",  6316 => x"4161003f",  6317 => x"31810020",
     6318 => x"78010001",  6319 => x"3821678c",  6320 => x"28230030",
     6321 => x"44600004",  6322 => x"b9600800",  6323 => x"b9801000",
     6324 => x"d8600000",  6325 => x"2b9d0004",  6326 => x"2b8b000c",
     6327 => x"2b8c0008",  6328 => x"379c000c",  6329 => x"c3a00000",
     6330 => x"2c230022",  6331 => x"0c430004",  6332 => x"28230024",
     6333 => x"58430000",  6334 => x"28210028",  6335 => x"58410008",
     6336 => x"c3a00000",  6337 => x"379cfff4",  6338 => x"5b8b000c",
     6339 => x"5b8c0008",  6340 => x"5b9d0004",  6341 => x"b8205800",
     6342 => x"2c210022",  6343 => x"b8406000",  6344 => x"34030008",
     6345 => x"0c410004",  6346 => x"29610024",  6347 => x"58410000",
     6348 => x"29610028",  6349 => x"58410008",  6350 => x"3441000c",
     6351 => x"3562002c",  6352 => x"f80032f3",  6353 => x"2d610034",
     6354 => x"0d810014",  6355 => x"2b9d0004",  6356 => x"2b8b000c",
     6357 => x"2b8c0008",  6358 => x"379c000c",  6359 => x"c3a00000",
     6360 => x"379cfff4",  6361 => x"5b8b000c",  6362 => x"5b8c0008",
     6363 => x"5b9d0004",  6364 => x"282b003c",  6365 => x"b8206000",
     6366 => x"34020000",  6367 => x"41610000",  6368 => x"3403000a",
     6369 => x"202100f0",  6370 => x"3821000b",  6371 => x"31610000",
     6372 => x"34010040",  6373 => x"0d610002",  6374 => x"2d810306",
     6375 => x"34210001",  6376 => x"2021ffff",  6377 => x"0d810306",
     6378 => x"0d61001e",  6379 => x"34010005",  6380 => x"31610020",
     6381 => x"298102c8",  6382 => x"4021000b",  6383 => x"31610021",
     6384 => x"35610022",  6385 => x"f8003350",  6386 => x"29810020",
     6387 => x"34030008",  6388 => x"28220018",  6389 => x"28210014",
     6390 => x"2c420000",  6391 => x"0d62002c",  6392 => x"4021001c",
     6393 => x"3161002f",  6394 => x"29810020",  6395 => x"28210014",
     6396 => x"40210018",  6397 => x"31610030",  6398 => x"29810020",
     6399 => x"28210014",  6400 => x"40210019",  6401 => x"31610031",
     6402 => x"29810020",  6403 => x"28210014",  6404 => x"2c22001a",
     6405 => x"0d620032",  6406 => x"4021001d",  6407 => x"31610034",
     6408 => x"29810020",  6409 => x"28220014",  6410 => x"35610035",
     6411 => x"34420010",  6412 => x"f80032b7",  6413 => x"29810020",
     6414 => x"28220010",  6415 => x"28210018",  6416 => x"2c420000",
     6417 => x"0d62003d",  6418 => x"4021001c",  6419 => x"34020040",
     6420 => x"3161003f",  6421 => x"78010001",  6422 => x"3821678c",
     6423 => x"2823002c",  6424 => x"44600004",  6425 => x"b9800800",
     6426 => x"d8600000",  6427 => x"b8201000",  6428 => x"b9800800",
     6429 => x"3403000b",  6430 => x"34040000",  6431 => x"fbfffebc",
     6432 => x"2b9d0004",  6433 => x"2b8b000c",  6434 => x"2b8c0008",
     6435 => x"379c000c",  6436 => x"c3a00000",  6437 => x"379cffc8",
     6438 => x"5b8b0018",  6439 => x"5b8c0014",  6440 => x"5b8d0010",
     6441 => x"5b8e000c",  6442 => x"5b8f0008",  6443 => x"5b9d0004",
     6444 => x"28220028",  6445 => x"378c001c",  6446 => x"b8205800",
     6447 => x"28430000",  6448 => x"b9801000",  6449 => x"378f0030",
     6450 => x"d8600000",  6451 => x"b9800800",  6452 => x"b9e01000",
     6453 => x"f8000103",  6454 => x"296c003c",  6455 => x"340efff0",
     6456 => x"340d002c",  6457 => x"41810000",  6458 => x"0d8d0002",
     6459 => x"34020000",  6460 => x"a02e0800",  6461 => x"31810000",
     6462 => x"2d6102f0",  6463 => x"34030008",  6464 => x"34210001",
     6465 => x"2021ffff",  6466 => x"0d6102f0",  6467 => x"31800020",
     6468 => x"0d81001e",  6469 => x"296102c8",  6470 => x"4021000d",
     6471 => x"31810021",  6472 => x"35810008",  6473 => x"f80032f8",
     6474 => x"2f810034",  6475 => x"3402002c",  6476 => x"34030000",
     6477 => x"0d810022",  6478 => x"2b810030",  6479 => x"34040001",
     6480 => x"59810024",  6481 => x"2b810038",  6482 => x"59810028",
     6483 => x"b9600800",  6484 => x"fbfffe87",  6485 => x"5c200023",
     6486 => x"29610020",  6487 => x"356c00f8",  6488 => x"b9801000",
     6489 => x"28230008",  6490 => x"b9800800",  6491 => x"34630018",
     6492 => x"f8000101",  6493 => x"b9e01000",  6494 => x"b9800800",
     6495 => x"f80000d9",  6496 => x"2961003c",  6497 => x"34030008",
     6498 => x"34040000",  6499 => x"40220000",  6500 => x"0c2d0002",
     6501 => x"a04e7000",  6502 => x"39ce0008",  6503 => x"302e0000",
     6504 => x"2d6202f0",  6505 => x"0c22001e",  6506 => x"34020002",
     6507 => x"30220020",  6508 => x"296202c8",  6509 => x"4042000d",
     6510 => x"30220021",  6511 => x"2f820034",  6512 => x"0c220022",
     6513 => x"2b820030",  6514 => x"58220024",  6515 => x"2b820038",
     6516 => x"58220028",  6517 => x"b9600800",  6518 => x"3402002c",
     6519 => x"fbfffe64",  6520 => x"2b9d0004",  6521 => x"2b8b0018",
     6522 => x"2b8c0014",  6523 => x"2b8d0010",  6524 => x"2b8e000c",
     6525 => x"2b8f0008",  6526 => x"379c0038",  6527 => x"c3a00000",
     6528 => x"379cffd4",  6529 => x"5b8b000c",  6530 => x"5b8c0008",
     6531 => x"5b9d0004",  6532 => x"28220028",  6533 => x"378b0010",
     6534 => x"b8206000",  6535 => x"28430000",  6536 => x"b9601000",
     6537 => x"d8600000",  6538 => x"37820024",  6539 => x"b9600800",
     6540 => x"f80000ac",  6541 => x"298b003c",  6542 => x"34020000",
     6543 => x"34030008",  6544 => x"41610000",  6545 => x"202100f0",
     6546 => x"38210001",  6547 => x"31610000",  6548 => x"3401002c",
     6549 => x"0d610002",  6550 => x"2d8102f2",  6551 => x"34210001",
     6552 => x"2021ffff",  6553 => x"0d8102f2",  6554 => x"0d61001e",
     6555 => x"34010001",  6556 => x"31610020",  6557 => x"3401007f",
     6558 => x"31610021",  6559 => x"35610008",  6560 => x"f80032a1",
     6561 => x"2f810028",  6562 => x"3402002c",  6563 => x"34030001",
     6564 => x"0d610022",  6565 => x"2b810024",  6566 => x"34040001",
     6567 => x"59610024",  6568 => x"2b81002c",  6569 => x"59610028",
     6570 => x"b9800800",  6571 => x"fbfffe30",  6572 => x"2b9d0004",
     6573 => x"2b8b000c",  6574 => x"2b8c0008",  6575 => x"379c002c",
     6576 => x"c3a00000",  6577 => x"379cffe8",  6578 => x"5b8b000c",
     6579 => x"5b8c0008",  6580 => x"5b9d0004",  6581 => x"b8206000",
     6582 => x"b8400800",  6583 => x"37820010",  6584 => x"f8000080",
     6585 => x"298b003c",  6586 => x"34020000",  6587 => x"34030008",
     6588 => x"41610000",  6589 => x"202100f0",  6590 => x"38210009",
     6591 => x"31610000",  6592 => x"34010036",  6593 => x"0d610002",
     6594 => x"41810312",  6595 => x"31610004",  6596 => x"35610008",
     6597 => x"f800327c",  6598 => x"2981031c",  6599 => x"35820320",
     6600 => x"34030008",  6601 => x"59610008",  6602 => x"29810318",
     6603 => x"5961000c",  6604 => x"2d81032a",  6605 => x"0d61001e",
     6606 => x"34010003",  6607 => x"31610020",  6608 => x"298102c8",
     6609 => x"4021000a",  6610 => x"31610021",  6611 => x"2f810014",
     6612 => x"0d610022",  6613 => x"2b810010",  6614 => x"59610024",
     6615 => x"2b810018",  6616 => x"59610028",  6617 => x"3561002c",
     6618 => x"f80031e9",  6619 => x"2d810328",  6620 => x"34020036",
     6621 => x"34030009",  6622 => x"0d610034",  6623 => x"34040000",
     6624 => x"b9800800",  6625 => x"fbfffdfa",  6626 => x"2b9d0004",
     6627 => x"2b8b000c",  6628 => x"2b8c0008",  6629 => x"379c0018",
     6630 => x"c3a00000",  6631 => x"379cfff0",  6632 => x"5b8b0010",
     6633 => x"5b8c000c",  6634 => x"5b8d0008",  6635 => x"5b9d0004",
     6636 => x"78030001",  6637 => x"282d0004",  6638 => x"38635a2c",
     6639 => x"28620000",  6640 => x"b8205800",  6641 => x"b9a00800",
     6642 => x"f8003123",  6643 => x"78030001",  6644 => x"296c0000",
     6645 => x"38635a2c",  6646 => x"28620000",  6647 => x"b42c6000",
     6648 => x"596c0000",  6649 => x"b9a00800",  6650 => x"f8003148",
     6651 => x"59610004",  6652 => x"4c0c0007",  6653 => x"4c20000f",
     6654 => x"358cffff",  6655 => x"78030001",  6656 => x"596c0000",
     6657 => x"38635a2c",  6658 => x"e0000007",  6659 => x"45800009",
     6660 => x"4c010008",  6661 => x"358c0001",  6662 => x"78030001",
     6663 => x"596c0000",  6664 => x"38635a40",  6665 => x"28620000",
     6666 => x"b4220800",  6667 => x"59610004",  6668 => x"2b9d0004",
     6669 => x"2b8b0010",  6670 => x"2b8c000c",  6671 => x"2b8d0008",
     6672 => x"379c0010",  6673 => x"c3a00000",  6674 => x"379cffe8",
     6675 => x"5b8b0008",  6676 => x"5b9d0004",  6677 => x"5b82000c",
     6678 => x"5b830010",  6679 => x"5b830014",  6680 => x"5b820018",
     6681 => x"b8205800",  6682 => x"4c600006",  6683 => x"78010001",
     6684 => x"78020001",  6685 => x"382145e4",  6686 => x"38425d20",
     6687 => x"f80017d0",  6688 => x"2b810018",  6689 => x"38028000",
     6690 => x"2b830014",  6691 => x"b4221000",  6692 => x"f4220800",
     6693 => x"00420010",  6694 => x"b4230800",  6695 => x"3c230010",
     6696 => x"00210010",  6697 => x"b8431000",  6698 => x"78030001",
     6699 => x"38635a2c",  6700 => x"5b820018",  6701 => x"28620000",
     6702 => x"5b810014",  6703 => x"37810014",  6704 => x"fbffec4a",
     6705 => x"59610004",  6706 => x"2b810018",  6707 => x"59610000",
     6708 => x"2b9d0004",  6709 => x"2b8b0008",  6710 => x"379c0018",
     6711 => x"c3a00000",  6712 => x"379cfffc",  6713 => x"5b9d0004",
     6714 => x"28230000",  6715 => x"48030003",  6716 => x"28210004",
     6717 => x"4c200006",  6718 => x"78010001",  6719 => x"38214610",
     6720 => x"f80017af",  6721 => x"3401ffff",  6722 => x"e0000005",
     6723 => x"58410008",  6724 => x"58430000",  6725 => x"0c400004",
     6726 => x"34010000",  6727 => x"2b9d0004",  6728 => x"379c0004",
     6729 => x"c3a00000",  6730 => x"379cfffc",  6731 => x"5b9d0004",
     6732 => x"78050001",  6733 => x"38a55a44",  6734 => x"28430000",
     6735 => x"28a40000",  6736 => x"54640006",  6737 => x"28420008",
     6738 => x"58230000",  6739 => x"58220004",  6740 => x"34010000",
     6741 => x"e0000005",  6742 => x"78010001",  6743 => x"3821464c",
     6744 => x"f8001797",  6745 => x"3401ffff",  6746 => x"2b9d0004",
     6747 => x"379c0004",  6748 => x"c3a00000",  6749 => x"379cfffc",
     6750 => x"5b9d0004",  6751 => x"28660000",  6752 => x"28450000",
     6753 => x"28630004",  6754 => x"28420004",  6755 => x"b4c52800",
     6756 => x"58250000",  6757 => x"b4621000",  6758 => x"58220004",
     6759 => x"fbffff80",  6760 => x"2b9d0004",  6761 => x"379c0004",
     6762 => x"c3a00000",  6763 => x"379cfffc",  6764 => x"5b9d0004",
     6765 => x"28460000",  6766 => x"28650000",  6767 => x"c8c52800",
     6768 => x"58250000",  6769 => x"28450004",  6770 => x"28620004",
     6771 => x"c8a21000",  6772 => x"58220004",  6773 => x"fbffff72",
     6774 => x"2b9d0004",  6775 => x"379c0004",  6776 => x"c3a00000",
     6777 => x"379cfffc",  6778 => x"5b9d0004",  6779 => x"78040001",
     6780 => x"38845a48",  6781 => x"28230000",  6782 => x"28820000",
     6783 => x"a0621000",  6784 => x"4c400005",  6785 => x"3442ffff",
     6786 => x"3404fffe",  6787 => x"b8441000",  6788 => x"34420001",
     6789 => x"78050001",  6790 => x"38a55a2c",  6791 => x"28a40000",
     6792 => x"88441000",  6793 => x"28240004",  6794 => x"b4441000",
     6795 => x"0064001f",  6796 => x"b4831800",  6797 => x"14630001",
     6798 => x"58230000",  6799 => x"0043001f",  6800 => x"b4621000",
     6801 => x"14420001",  6802 => x"58220004",  6803 => x"fbffff54",
     6804 => x"2b9d0004",  6805 => x"379c0004",  6806 => x"c3a00000",
     6807 => x"379cfff8",  6808 => x"5b8b0008",  6809 => x"5b9d0004",
     6810 => x"28250000",  6811 => x"78030001",  6812 => x"b8201000",
     6813 => x"3863469c",  6814 => x"4805000a",  6815 => x"78030001",
     6816 => x"38634e44",  6817 => x"5ca00007",  6818 => x"28210004",
     6819 => x"78030001",  6820 => x"3863469c",  6821 => x"48a10003",
     6822 => x"78030001",  6823 => x"38634e44",  6824 => x"28410004",
     6825 => x"14a4001f",  6826 => x"780b0001",  6827 => x"1426001f",
     6828 => x"98853800",  6829 => x"396b7a88",  6830 => x"98c12800",
     6831 => x"78020001",  6832 => x"b9600800",  6833 => x"384246a0",
     6834 => x"c8e42000",  6835 => x"c8a62800",  6836 => x"f800172d",
     6837 => x"b9600800",  6838 => x"2b9d0004",  6839 => x"2b8b0008",
     6840 => x"379c0008",  6841 => x"c3a00000",  6842 => x"379cfff8",
     6843 => x"5b8b0008",  6844 => x"5b9d0004",  6845 => x"28220020",
     6846 => x"28240028",  6847 => x"b8205800",  6848 => x"28430004",
     6849 => x"58600038",  6850 => x"28430014",  6851 => x"0c20010c",
     6852 => x"0c600008",  6853 => x"28830014",  6854 => x"44600013",
     6855 => x"d8600000",  6856 => x"3402ffff",  6857 => x"5c220008",
     6858 => x"78040001",  6859 => x"b9600800",  6860 => x"34020004",
     6861 => x"34030001",  6862 => x"388446ac",  6863 => x"fbffe783",
     6864 => x"34010000",  6865 => x"29620020",  6866 => x"c8010800",
     6867 => x"3c21000a",  6868 => x"28420004",  6869 => x"1423001f",
     6870 => x"5841002c",  6871 => x"58430028",  6872 => x"e000000d",
     6873 => x"28420008",  6874 => x"28420038",  6875 => x"20420001",
     6876 => x"5c430005",  6877 => x"28840008",  6878 => x"34020000",
     6879 => x"34030000",  6880 => x"d8800000",  6881 => x"29610020",
     6882 => x"28210004",  6883 => x"58200028",  6884 => x"5820002c",
     6885 => x"29610020",  6886 => x"78040001",  6887 => x"34020004",
     6888 => x"28260004",  6889 => x"34030001",  6890 => x"b9600800",
     6891 => x"28c50028",  6892 => x"28c6002c",  6893 => x"388446c8",
     6894 => x"fbffe764",  6895 => x"2b9d0004",  6896 => x"2b8b0008",
     6897 => x"379c0008",  6898 => x"c3a00000",  6899 => x"379cfff0",
     6900 => x"5b8b0010",  6901 => x"5b8c000c",  6902 => x"5b8d0008",
     6903 => x"5b9d0004",  6904 => x"b8205800",  6905 => x"28210020",
     6906 => x"35620094",  6907 => x"35630080",  6908 => x"282d0004",
     6909 => x"356c00d0",  6910 => x"b9a00800",  6911 => x"fbffff6c",
     6912 => x"b9a01000",  6913 => x"b9801800",  6914 => x"b9a00800",
     6915 => x"fbffff68",  6916 => x"b9800800",  6917 => x"fbffff92",
     6918 => x"78040001",  6919 => x"b8202800",  6920 => x"34020004",
     6921 => x"b9600800",  6922 => x"34030003",  6923 => x"388446e8",
     6924 => x"fbffe746",  6925 => x"2b9d0004",  6926 => x"2b8b0010",
     6927 => x"2b8c000c",  6928 => x"2b8d0008",  6929 => x"379c0010",
     6930 => x"c3a00000",  6931 => x"379cffb8",  6932 => x"5b8b0024",
     6933 => x"5b8c0020",  6934 => x"5b8d001c",  6935 => x"5b8e0018",
     6936 => x"5b8f0014",  6937 => x"5b900010",  6938 => x"5b91000c",
     6939 => x"5b920008",  6940 => x"5b9d0004",  6941 => x"28220020",
     6942 => x"b8205800",  6943 => x"284d0004",  6944 => x"284c0010",
     6945 => x"28220080",  6946 => x"5c400008",  6947 => x"28230084",
     6948 => x"5c620006",  6949 => x"78040001",  6950 => x"34020004",
     6951 => x"34030002",  6952 => x"38844700",  6953 => x"e000006e",
     6954 => x"35af0014",  6955 => x"357000bc",  6956 => x"357100a8",
     6957 => x"b9e00800",  6958 => x"ba001000",  6959 => x"ba201800",
     6960 => x"fbffff3b",  6961 => x"357200d0",  6962 => x"b9e01000",
     6963 => x"ba401800",  6964 => x"b9e00800",  6965 => x"fbffff36",
     6966 => x"ba400800",  6967 => x"fbffff60",  6968 => x"78040001",
     6969 => x"b8202800",  6970 => x"34020004",  6971 => x"34030003",
     6972 => x"38844720",  6973 => x"b9600800",  6974 => x"fbffe714",
     6975 => x"35610080",  6976 => x"fbffff57",  6977 => x"78040001",
     6978 => x"b8202800",  6979 => x"34020004",  6980 => x"34030002",
     6981 => x"38844738",  6982 => x"b9600800",  6983 => x"fbffe70b",
     6984 => x"35610094",  6985 => x"fbffff4e",  6986 => x"78040001",
     6987 => x"b8202800",  6988 => x"34020004",  6989 => x"34030002",
     6990 => x"38844740",  6991 => x"b9600800",  6992 => x"fbffe702",
     6993 => x"ba200800",  6994 => x"fbffff45",  6995 => x"78040001",
     6996 => x"b8202800",  6997 => x"34020004",  6998 => x"34030002",
     6999 => x"38844748",  7000 => x"b9600800",  7001 => x"fbffe6f9",
     7002 => x"ba000800",  7003 => x"fbffff3c",  7004 => x"78040001",
     7005 => x"b8202800",  7006 => x"34020004",  7007 => x"34030002",
     7008 => x"38844750",  7009 => x"b9600800",  7010 => x"fbffe6f0",
     7011 => x"b9a00800",  7012 => x"fbffff33",  7013 => x"78040001",
     7014 => x"b8202800",  7015 => x"34020004",  7016 => x"34030001",
     7017 => x"38844758",  7018 => x"b9600800",  7019 => x"fbffe6e7",
     7020 => x"b9e00800",  7021 => x"fbffff2a",  7022 => x"78040001",
     7023 => x"b8202800",  7024 => x"38844770",  7025 => x"b9600800",
     7026 => x"34020004",  7027 => x"34030001",  7028 => x"fbffe6de",
     7029 => x"29610020",  7030 => x"358e0018",  7031 => x"28220004",
     7032 => x"b9c00800",  7033 => x"34430014",  7034 => x"fbfffee3",
     7035 => x"b9c00800",  7036 => x"fbfffefd",  7037 => x"b9c00800",
     7038 => x"fbffff19",  7039 => x"78040001",  7040 => x"b8202800",
     7041 => x"34020004",  7042 => x"b9600800",  7043 => x"34030001",
     7044 => x"38844788",  7045 => x"fbffe6cd",  7046 => x"29610020",
     7047 => x"28220010",  7048 => x"28260004",  7049 => x"28420018",
     7050 => x"5c400142",  7051 => x"28210008",  7052 => x"28270030",
     7053 => x"44e2013c",  7054 => x"28c20000",  7055 => x"5c400003",
     7056 => x"28c30014",  7057 => x"44620008",  7058 => x"78040001",
     7059 => x"b9600800",  7060 => x"34020004",  7061 => x"34030001",
     7062 => x"3884479c",  7063 => x"fbffe6bb",  7064 => x"e0000134",
     7065 => x"28c50004",  7066 => x"48a70003",  7067 => x"28c20018",
     7068 => x"4ce2012d",  7069 => x"28c60018",  7070 => x"78040001",
     7071 => x"b9600800",  7072 => x"34020004",  7073 => x"34030001",
     7074 => x"388447c8",  7075 => x"fbffe6af",  7076 => x"e0000128",
     7077 => x"2982001c",  7078 => x"59a20034",  7079 => x"1c220040",
     7080 => x"29a10034",  7081 => x"3444ffff",  7082 => x"1423001f",
     7083 => x"98612800",  7084 => x"c8a32800",  7085 => x"3403001f",
     7086 => x"c8621800",  7087 => x"94a33800",  7088 => x"34820001",
     7089 => x"34630001",  7090 => x"3484ffff",  7091 => x"5ce0fffc",
     7092 => x"34030001",  7093 => x"bc621000",  7094 => x"4c460002",
     7095 => x"59a20038",  7096 => x"29a30038",  7097 => x"4c620003",
     7098 => x"34630001",  7099 => x"59a30038",  7100 => x"2982001c",
     7101 => x"4c400002",  7102 => x"5981001c",  7103 => x"2982001c",
     7104 => x"4c400002",  7105 => x"5980001c",  7106 => x"2985001c",
     7107 => x"08210003",  7108 => x"4c25000d",  7109 => x"78040001",
     7110 => x"b9600800",  7111 => x"34020004",  7112 => x"34030001",
     7113 => x"3884480c",  7114 => x"fbffe688",  7115 => x"29a10034",
     7116 => x"29a20038",  7117 => x"3c210001",  7118 => x"34420001",
     7119 => x"b4410800",  7120 => x"5981001c",  7121 => x"29af0038",
     7122 => x"29a20034",  7123 => x"35900004",  7124 => x"35e1ffff",
     7125 => x"88220800",  7126 => x"2982001c",  7127 => x"b4220800",
     7128 => x"b9e01000",  7129 => x"f8002f3c",  7130 => x"59a10034",
     7131 => x"78040001",  7132 => x"b8203000",  7133 => x"b9e02800",
     7134 => x"38844824",  7135 => x"5981001c",  7136 => x"34020004",
     7137 => x"b9600800",  7138 => x"34030001",  7139 => x"fbffe66f",
     7140 => x"b9a01000",  7141 => x"b9c01800",  7142 => x"ba000800",
     7143 => x"fbfffe84",  7144 => x"ba000800",  7145 => x"fbfffeae",
     7146 => x"78040001",  7147 => x"b8202800",  7148 => x"34020004",
     7149 => x"b9600800",  7150 => x"34030001",  7151 => x"38844848",
     7152 => x"fbffe662",  7153 => x"296f0020",  7154 => x"29e10008",
     7155 => x"2825002c",  7156 => x"44a00011",  7157 => x"29820004",
     7158 => x"44400007",  7159 => x"78040001",  7160 => x"b9600800",
     7161 => x"34020004",  7162 => x"34030001",  7163 => x"38844864",
     7164 => x"e3ffff9b",  7165 => x"29820008",  7166 => x"4ca20007",
     7167 => x"78040001",  7168 => x"b9600800",  7169 => x"34020004",
     7170 => x"34030001",  7171 => x"38844894",  7172 => x"e00000c3",
     7173 => x"29820004",  7174 => x"44400031",  7175 => x"28220038",
     7176 => x"20410001",  7177 => x"5c2000c3",  7178 => x"20420002",
     7179 => x"5c410019",  7180 => x"296300c4",  7181 => x"296200c8",
     7182 => x"296100cc",  7183 => x"5b830030",  7184 => x"29e30010",
     7185 => x"296500bc",  7186 => x"296400c0",  7187 => x"378c0028",
     7188 => x"5b820034",  7189 => x"5b810038",  7190 => x"b9801000",
     7191 => x"b9800800",  7192 => x"34630018",  7193 => x"5b850028",
     7194 => x"5b84002c",  7195 => x"fbfffe42",  7196 => x"29610028",
     7197 => x"b9801000",  7198 => x"28230004",  7199 => x"b9600800",
     7200 => x"d8600000",  7201 => x"b9600800",  7202 => x"fbfffe98",
     7203 => x"e00000a9",  7204 => x"29820008",  7205 => x"78030001",
     7206 => x"38635a4c",  7207 => x"28610000",  7208 => x"ec021000",
     7209 => x"78050001",  7210 => x"c8021000",  7211 => x"38a55a50",
     7212 => x"a0411000",  7213 => x"28a10000",  7214 => x"b4411000",
     7215 => x"29610028",  7216 => x"c8021000",  7217 => x"28230010",
     7218 => x"5c600002",  7219 => x"2823000c",  7220 => x"b9600800",
     7221 => x"d8600000",  7222 => x"e0000096",  7223 => x"29830008",
     7224 => x"29ed0004",  7225 => x"78050001",  7226 => x"1462001f",
     7227 => x"29b0002c",  7228 => x"00640016",  7229 => x"3c63000a",
     7230 => x"29ae0028",  7231 => x"3c42000a",  7232 => x"b4708000",
     7233 => x"b8821000",  7234 => x"f4701800",  7235 => x"b44e1000",
     7236 => x"b4627000",  7237 => x"1c22003e",  7238 => x"38a55a50",
     7239 => x"28a40000",  7240 => x"1441001f",  7241 => x"34030000",
     7242 => x"59ae0028",  7243 => x"59b0002c",  7244 => x"f8002ea2",
     7245 => x"00430016",  7246 => x"3c21000a",  7247 => x"3c42000a",
     7248 => x"b8610800",  7249 => x"49c1000b",  7250 => x"5dc10002",
     7251 => x"56020009",  7252 => x"c8021000",  7253 => x"7c430000",
     7254 => x"c8010800",  7255 => x"c8230800",  7256 => x"482e0004",
     7257 => x"5c2e0005",  7258 => x"54500002",  7259 => x"e0000003",
     7260 => x"59a10028",  7261 => x"59a2002c",  7262 => x"29a10028",
     7263 => x"29a2002c",  7264 => x"48200003",  7265 => x"5c200004",
     7266 => x"44410003",  7267 => x"340d0000",  7268 => x"e0000002",
     7269 => x"340dffff",  7270 => x"5b810044",  7271 => x"5b820048",
     7272 => x"45a00007",  7273 => x"c8021000",  7274 => x"7c430000",
     7275 => x"c8010800",  7276 => x"c8230800",  7277 => x"5b810044",
     7278 => x"5b820048",  7279 => x"29e20008",  7280 => x"37810044",
     7281 => x"1c42003e",  7282 => x"fbffea08",  7283 => x"45a00009",
     7284 => x"2b810048",  7285 => x"2b820044",  7286 => x"c8010800",
     7287 => x"7c230000",  7288 => x"c8021000",  7289 => x"c8431000",
     7290 => x"5b820044",  7291 => x"5b810048",  7292 => x"29820008",
     7293 => x"1441001f",  7294 => x"00430016",  7295 => x"3c21000a",
     7296 => x"ec026000",  7297 => x"3c42000a",  7298 => x"b8610800",
     7299 => x"c80c6000",  7300 => x"5b81003c",  7301 => x"5b820040",
     7302 => x"45800007",  7303 => x"c8021000",  7304 => x"7c430000",
     7305 => x"c8010800",  7306 => x"c8230800",  7307 => x"5b81003c",
     7308 => x"5b820040",  7309 => x"29610020",  7310 => x"28220008",
     7311 => x"3781003c",  7312 => x"1c42003c",  7313 => x"fbffe9e9",
     7314 => x"45800009",  7315 => x"2b810040",  7316 => x"2b82003c",
     7317 => x"c8010800",  7318 => x"7c230000",  7319 => x"c8021000",
     7320 => x"c8431000",  7321 => x"5b82003c",  7322 => x"5b810040",
     7323 => x"2b830048",  7324 => x"2b820040",  7325 => x"2b81003c",
     7326 => x"2b840044",  7327 => x"b4621000",  7328 => x"f4621800",
     7329 => x"b4810800",  7330 => x"b4610800",  7331 => x"48200003",
     7332 => x"5c200006",  7333 => x"44410005",  7334 => x"3c210016",
     7335 => x"0042000a",  7336 => x"b8221000",  7337 => x"e0000009",
     7338 => x"c8021000",  7339 => x"7c430000",  7340 => x"c8010800",
     7341 => x"c8230800",  7342 => x"3c210016",  7343 => x"0042000a",
     7344 => x"b8221000",  7345 => x"c8021000",  7346 => x"29610020",
     7347 => x"28210008",  7348 => x"28250038",  7349 => x"20a50001",
     7350 => x"5ca00008",  7351 => x"29640028",  7352 => x"c8021000",
     7353 => x"28830010",  7354 => x"5c650002",  7355 => x"2883000c",
     7356 => x"b9600800",  7357 => x"d8600000",  7358 => x"29610020",
     7359 => x"78040001",  7360 => x"34020004",  7361 => x"28210004",
     7362 => x"34030002",  7363 => x"388448d0",  7364 => x"2825002c",
     7365 => x"b9600800",  7366 => x"14a5000a",  7367 => x"fbffe58b",
     7368 => x"e0000004",  7369 => x"29a60038",  7370 => x"4c06fedb",
     7371 => x"e3fffedc",  7372 => x"2b9d0004",  7373 => x"2b8b0024",
     7374 => x"2b8c0020",  7375 => x"2b8d001c",  7376 => x"2b8e0018",
     7377 => x"2b8f0014",  7378 => x"2b900010",  7379 => x"2b91000c",
     7380 => x"2b920008",  7381 => x"379c0048",  7382 => x"c3a00000",
     7383 => x"379cfffc",  7384 => x"5b9d0004",  7385 => x"78030001",
     7386 => x"3c420002",  7387 => x"38636804",  7388 => x"b4622800",
     7389 => x"28a50000",  7390 => x"78040001",  7391 => x"34020006",
     7392 => x"34030001",  7393 => x"388448e8",  7394 => x"fbffe570",
     7395 => x"2b9d0004",  7396 => x"379c0004",  7397 => x"c3a00000",
     7398 => x"379cfff0",  7399 => x"5b8b0010",  7400 => x"5b8c000c",
     7401 => x"5b8d0008",  7402 => x"5b9d0004",  7403 => x"b8205800",
     7404 => x"78010001",  7405 => x"38217aa0",  7406 => x"b8406800",
     7407 => x"28220000",  7408 => x"5c400005",  7409 => x"29620020",
     7410 => x"2844000c",  7411 => x"28820008",  7412 => x"58220000",
     7413 => x"78040001",  7414 => x"78010001",  7415 => x"38847aa0",
     7416 => x"38215a54",  7417 => x"28260000",  7418 => x"28850000",
     7419 => x"340c0190",  7420 => x"bd836000",  7421 => x"88a62800",
     7422 => x"b9801000",  7423 => x"34a53039",  7424 => x"00a10010",
     7425 => x"88a62800",  7426 => x"202107ff",  7427 => x"34a53039",
     7428 => x"58850000",  7429 => x"00a50010",  7430 => x"3c24000a",
     7431 => x"20a103ff",  7432 => x"b8240800",  7433 => x"f8002e69",
     7434 => x"3d820001",  7435 => x"b4221000",  7436 => x"29610028",
     7437 => x"28230018",  7438 => x"b9600800",  7439 => x"d8600000",
     7440 => x"35a200b2",  7441 => x"3c420002",  7442 => x"b5625800",
     7443 => x"59610004",  7444 => x"2b9d0004",  7445 => x"2b8b0010",
     7446 => x"2b8c000c",  7447 => x"2b8d0008",  7448 => x"379c0010",
     7449 => x"c3a00000",  7450 => x"379cfff0",  7451 => x"5b8b0010",
     7452 => x"5b8c000c",  7453 => x"5b8d0008",  7454 => x"5b9d0004",
     7455 => x"282b000c",  7456 => x"b8206000",  7457 => x"34010001",
     7458 => x"59610000",  7459 => x"29810024",  7460 => x"48200002",
     7461 => x"34010001",  7462 => x"0d61000c",  7463 => x"29810008",
     7464 => x"5c200002",  7465 => x"59820008",  7466 => x"298d0008",
     7467 => x"3561000e",  7468 => x"34030004",  7469 => x"b9a01000",
     7470 => x"f8002e95",  7471 => x"2d62000c",  7472 => x"34010001",
     7473 => x"5c410004",  7474 => x"29810000",  7475 => x"4021001d",
     7476 => x"64210002",  7477 => x"59610018",  7478 => x"41a10044",
     7479 => x"2d67000c",  7480 => x"34060002",  7481 => x"31610012",
     7482 => x"41a10045",  7483 => x"34050001",  7484 => x"3404ffff",
     7485 => x"31610013",  7486 => x"41a10046",  7487 => x"31610014",
     7488 => x"34010000",  7489 => x"e000000c",  7490 => x"08220374",
     7491 => x"29880000",  7492 => x"b5021000",  7493 => x"44600004",
     7494 => x"4043001d",  7495 => x"44660002",  7496 => x"59600018",
     7497 => x"58410338",  7498 => x"58450000",  7499 => x"0c44010e",
     7500 => x"34210001",  7501 => x"29630018",  7502 => x"48e1fff4",
     7503 => x"44600006",  7504 => x"78010001",  7505 => x"38214978",
     7506 => x"f800149d",  7507 => x"3401ffff",  7508 => x"3161000e",
     7509 => x"78010001",  7510 => x"3821678c",  7511 => x"28230004",
     7512 => x"34010000",  7513 => x"44600004",  7514 => x"b9800800",
     7515 => x"b9a01000",  7516 => x"d8600000",  7517 => x"2b9d0004",
     7518 => x"2b8b0010",  7519 => x"2b8c000c",  7520 => x"2b8d0008",
     7521 => x"379c0010",  7522 => x"c3a00000",  7523 => x"379cfffc",
     7524 => x"5b9d0004",  7525 => x"78020001",  7526 => x"3842678c",
     7527 => x"28430008",  7528 => x"34020000",  7529 => x"44600003",
     7530 => x"d8600000",  7531 => x"b8201000",  7532 => x"b8400800",
     7533 => x"2b9d0004",  7534 => x"379c0004",  7535 => x"c3a00000",
     7536 => x"78010001",  7537 => x"38216870",  7538 => x"28220000",
     7539 => x"78010001",  7540 => x"38216654",  7541 => x"e0000004",
     7542 => x"28440000",  7543 => x"44640004",  7544 => x"3421000c",
     7545 => x"28230000",  7546 => x"5c60fffc",  7547 => x"28210004",
     7548 => x"c3a00000",  7549 => x"379cfff4",  7550 => x"5b9d0004",
     7551 => x"5b810008",  7552 => x"5b82000c",  7553 => x"b8401800",
     7554 => x"5c20000b",  7555 => x"78020001",  7556 => x"38425a3c",
     7557 => x"28410000",  7558 => x"54610007",  7559 => x"78010001",
     7560 => x"78020001",  7561 => x"3842499c",  7562 => x"38217aa8",
     7563 => x"f8001456",  7564 => x"e000000d",  7565 => x"78030001",
     7566 => x"38635a2c",  7567 => x"28620000",  7568 => x"37810008",
     7569 => x"fbffe8e9",  7570 => x"2b83000c",  7571 => x"b8202000",
     7572 => x"78020001",  7573 => x"78010001",  7574 => x"38217aa8",
     7575 => x"384249a0",  7576 => x"f8001449",  7577 => x"78010001",
     7578 => x"38217aa8",  7579 => x"2b9d0004",  7580 => x"379c000c",
     7581 => x"c3a00000",  7582 => x"379cff18",  7583 => x"5b8b000c",
     7584 => x"5b8c0008",  7585 => x"5b9d0004",  7586 => x"78010001",
     7587 => x"38216870",  7588 => x"28210000",  7589 => x"282b0014",
     7590 => x"78010001",  7591 => x"38219290",  7592 => x"28220000",
     7593 => x"34010000",  7594 => x"444000ce",  7595 => x"780c0001",
     7596 => x"398c7aa4",  7597 => x"29810000",  7598 => x"5c200008",
     7599 => x"f8001a00",  7600 => x"78020001",  7601 => x"38426168",
     7602 => x"28420000",  7603 => x"a4401000",  7604 => x"b4410800",
     7605 => x"59810000",  7606 => x"78010001",  7607 => x"38218f2c",
     7608 => x"28210000",  7609 => x"296200b8",  7610 => x"5c220007",
     7611 => x"78010001",  7612 => x"38217594",  7613 => x"28230000",
     7614 => x"34020003",  7615 => x"34010000",  7616 => x"446200b8",
     7617 => x"f80019ee",  7618 => x"78030001",  7619 => x"78020001",
     7620 => x"38636168",  7621 => x"38427aa4",  7622 => x"28630000",
     7623 => x"28420000",  7624 => x"b4621000",  7625 => x"c8220800",
     7626 => x"4c200007",  7627 => x"78010001",  7628 => x"38217594",
     7629 => x"28230000",  7630 => x"34020003",  7631 => x"34010000",
     7632 => x"5c6200a8",  7633 => x"f80019de",  7634 => x"78020001",
     7635 => x"38427aa4",  7636 => x"58410000",  7637 => x"296200b8",
     7638 => x"78010001",  7639 => x"38218f2c",  7640 => x"58220000",
     7641 => x"378100d8",  7642 => x"378200e0",  7643 => x"f8001d70",
     7644 => x"34020000",  7645 => x"37810010",  7646 => x"f8000287",
     7647 => x"378100e8",  7648 => x"378200e4",  7649 => x"f80019b5",
     7650 => x"2b8300e4",  7651 => x"2b8400e8",  7652 => x"2b82003c",
     7653 => x"78010001",  7654 => x"382149a8",  7655 => x"f8001408",
     7656 => x"2b820044",  7657 => x"78010001",  7658 => x"382149bc",
     7659 => x"7c420000",  7660 => x"f8001403",  7661 => x"fbffff83",
     7662 => x"b8201000",  7663 => x"78010001",  7664 => x"382149c8",
     7665 => x"f80013fe",  7666 => x"78010001",  7667 => x"38217594",
     7668 => x"28220000",  7669 => x"34010003",  7670 => x"5c41000a",
     7671 => x"29620010",  7672 => x"78010001",  7673 => x"382149d0",
     7674 => x"20420001",  7675 => x"f80013f4",  7676 => x"78010001",
     7677 => x"382149d8",  7678 => x"356200c0",  7679 => x"f80013f0",
     7680 => x"34010000",  7681 => x"f8002ae0",  7682 => x"b8201000",
     7683 => x"78010001",  7684 => x"382149e4",  7685 => x"f80013ea",
     7686 => x"2b8200dc",  7687 => x"2b8300e0",  7688 => x"78010001",
     7689 => x"382149ec",  7690 => x"f80013e5",  7691 => x"78010001",
     7692 => x"38217594",  7693 => x"28220000",  7694 => x"34010003",
     7695 => x"5c41004b",  7696 => x"296200a4",  7697 => x"296100a0",
     7698 => x"fbffff6b",  7699 => x"b8201000",  7700 => x"78010001",
     7701 => x"382149fc",  7702 => x"f80013d9",  7703 => x"296200b4",
     7704 => x"296100b0",  7705 => x"fbffff64",  7706 => x"b8201000",
     7707 => x"78010001",  7708 => x"38214a04",  7709 => x"f80013d2",
     7710 => x"29620018",  7711 => x"2963001c",  7712 => x"78010001",
     7713 => x"38214a0c",  7714 => x"f80013cd",  7715 => x"29620020",
     7716 => x"29630024",  7717 => x"78010001",  7718 => x"38214a20",
     7719 => x"f80013c8",  7720 => x"296200b4",  7721 => x"296300a4",
     7722 => x"78010001",  7723 => x"3c420001",  7724 => x"38214a34",
     7725 => x"c8621000",  7726 => x"f80013c1",  7727 => x"29620018",
     7728 => x"296100a4",  7729 => x"296300a0",  7730 => x"1444001f",
     7731 => x"c8221000",  7732 => x"f4410800",  7733 => x"c8641800",
     7734 => x"c8611800",  7735 => x"2961001c",  7736 => x"1424001f",
     7737 => x"c8410800",  7738 => x"f4221000",  7739 => x"c8641800",
     7740 => x"c8621000",  7741 => x"29630020",  7742 => x"1464001f",
     7743 => x"c8231800",  7744 => x"f4610800",  7745 => x"c8441000",
     7746 => x"c8410800",  7747 => x"29620024",  7748 => x"1444001f",
     7749 => x"c8621000",  7750 => x"f4431800",  7751 => x"c8240800",
     7752 => x"c8230800",  7753 => x"fbffff34",  7754 => x"b8201000",
     7755 => x"78010001",  7756 => x"38214a40",  7757 => x"f80013a2",
     7758 => x"296200ec",  7759 => x"78010001",  7760 => x"38214a4c",
     7761 => x"f800139e",  7762 => x"296200a8",  7763 => x"78010001",
     7764 => x"38214a54",  7765 => x"f800139a",  7766 => x"296200b8",
     7767 => x"78010001",  7768 => x"38214a60",  7769 => x"f8001396",
     7770 => x"3401ffff",  7771 => x"f8002a91",  7772 => x"b8206000",
     7773 => x"34010000",  7774 => x"f8002a8e",  7775 => x"b8205800",
     7776 => x"34010001",  7777 => x"f8002a8b",  7778 => x"78050001",
     7779 => x"b8202000",  7780 => x"b8a00800",  7781 => x"b9801000",
     7782 => x"b9601800",  7783 => x"38214a6c",  7784 => x"f8001387",
     7785 => x"78010001",  7786 => x"38214a80",  7787 => x"f8001bdb",
     7788 => x"2023ffff",  7789 => x"08632710",  7790 => x"b8201000",
     7791 => x"14420010",  7792 => x"14630010",  7793 => x"78010001",
     7794 => x"38214a84",  7795 => x"f800137c",  7796 => x"78010001",
     7797 => x"38214d20",  7798 => x"f8001379",  7799 => x"34010001",
     7800 => x"2b9d0004",  7801 => x"2b8b000c",  7802 => x"2b8c0008",
     7803 => x"379c00e8",  7804 => x"c3a00000",  7805 => x"379cfff4",
     7806 => x"5b8b000c",  7807 => x"5b8c0008",  7808 => x"5b9d0004",
     7809 => x"780b0001",  7810 => x"396b6870",  7811 => x"29610000",
     7812 => x"78020001",  7813 => x"38424a94",  7814 => x"282c0014",
     7815 => x"34010004",  7816 => x"f8000938",  7817 => x"fbfffee7",
     7818 => x"78020001",  7819 => x"b8201800",  7820 => x"38424aa4",
     7821 => x"34010007",  7822 => x"f8000932",  7823 => x"29810010",
     7824 => x"44200005",  7825 => x"29610000",  7826 => x"28220000",
     7827 => x"34010009",  7828 => x"44410007",  7829 => x"78020001",
     7830 => x"34010001",  7831 => x"38424aa8",  7832 => x"f8000928",
     7833 => x"34010000",  7834 => x"e0000006",  7835 => x"78020001",
     7836 => x"34010004",  7837 => x"38424ac0",  7838 => x"f8000922",
     7839 => x"34010001",  7840 => x"2b9d0004",  7841 => x"2b8b000c",
     7842 => x"2b8c0008",  7843 => x"379c000c",  7844 => x"c3a00000",
     7845 => x"379cfef0",  7846 => x"5b8b0018",  7847 => x"5b8c0014",
     7848 => x"5b8d0010",  7849 => x"5b8e000c",  7850 => x"5b8f0008",
     7851 => x"5b9d0004",  7852 => x"78010001",  7853 => x"38216870",
     7854 => x"28210000",  7855 => x"780c0001",  7856 => x"398c7ac4",
     7857 => x"282b0014",  7858 => x"29810000",  7859 => x"5c200008",
     7860 => x"f80018fb",  7861 => x"78020001",  7862 => x"38426168",
     7863 => x"28420000",  7864 => x"a4401000",  7865 => x"b4410800",
     7866 => x"59810000",  7867 => x"f80018f4",  7868 => x"78030001",
     7869 => x"78020001",  7870 => x"38636168",  7871 => x"38427ac4",
     7872 => x"28630000",  7873 => x"28420000",  7874 => x"b4621000",
     7875 => x"c8220800",  7876 => x"4c200007",  7877 => x"78010001",
     7878 => x"38217ac0",  7879 => x"28210000",  7880 => x"296200b8",
     7881 => x"340d0000",  7882 => x"44220192",  7883 => x"f80018e4",
     7884 => x"78020001",  7885 => x"38427ac4",  7886 => x"58410000",
     7887 => x"296200b8",  7888 => x"78010001",  7889 => x"38217ac0",
     7890 => x"58220000",  7891 => x"f8000933",  7892 => x"78040001",
     7893 => x"34010001",  7894 => x"34020001",  7895 => x"34030004",
     7896 => x"38844adc",  7897 => x"f8000906",  7898 => x"78040001",
     7899 => x"38844afc",  7900 => x"34030087",  7901 => x"34010002",
     7902 => x"34020001",  7903 => x"f8000900",  7904 => x"378100fc",
     7905 => x"37820108",  7906 => x"f8001c69",  7907 => x"78020001",
     7908 => x"34010004",  7909 => x"38424b08",  7910 => x"f80008da",
     7911 => x"2b820100",  7912 => x"2b8100fc",  7913 => x"34030000",
     7914 => x"f8000825",  7915 => x"78020001",  7916 => x"b8201800",
     7917 => x"38424aa4",  7918 => x"34010007",  7919 => x"f80008d1",
     7920 => x"34020000",  7921 => x"37810020",  7922 => x"f8000173",
     7923 => x"78040001",  7924 => x"34010004",  7925 => x"34020001",
     7926 => x"34030004",  7927 => x"38844b28",  7928 => x"f80008e7",
     7929 => x"78040001",  7930 => x"78050001",  7931 => x"34010006",
     7932 => x"34020001",  7933 => x"34030007",  7934 => x"38844b38",
     7935 => x"38a54b40",  7936 => x"f80008df",  7937 => x"2b81004c",
     7938 => x"44200005",  7939 => x"78020001",  7940 => x"34010002",
     7941 => x"38424b48",  7942 => x"e0000004",  7943 => x"78020001",
     7944 => x"34010001",  7945 => x"38424b54",  7946 => x"f80008b6",
     7947 => x"2b81004c",  7948 => x"4420014c",  7949 => x"37810110",
     7950 => x"3782010c",  7951 => x"f8001887",  7952 => x"2b83010c",
     7953 => x"2b840110",  7954 => x"78020001",  7955 => x"34010087",
     7956 => x"38424b60",  7957 => x"780c0001",  7958 => x"f80008aa",
     7959 => x"398c6870",  7960 => x"29810000",  7961 => x"282102c8",
     7962 => x"28210010",  7963 => x"282e0008",  7964 => x"5dc00039",
     7965 => x"78020001",  7966 => x"34010001",  7967 => x"38424b7c",
     7968 => x"f80008a0",  7969 => x"fbffff5c",  7970 => x"340d0001",
     7971 => x"442e0139",  7972 => x"78020001",  7973 => x"34010087",
     7974 => x"38424b84",  7975 => x"f8000899",  7976 => x"29810000",
     7977 => x"28210020",  7978 => x"28240010",  7979 => x"28830004",
     7980 => x"4460000b",  7981 => x"78020001",  7982 => x"38424ba4",
     7983 => x"28840008",  7984 => x"4c030003",  7985 => x"34010007",
     7986 => x"e0000003",  7987 => x"34010007",  7988 => x"c8042000",
     7989 => x"f800088b",  7990 => x"e0000126",  7991 => x"28830008",
     7992 => x"780b0001",  7993 => x"396b4bb0",  7994 => x"b9601000",
     7995 => x"34010007",  7996 => x"f8000884",  7997 => x"78020001",
     7998 => x"34010087",  7999 => x"38424bb8",  8000 => x"f8000880",
     8001 => x"29810000",  8002 => x"b9601000",  8003 => x"28210020",
     8004 => x"28230010",  8005 => x"34010007",  8006 => x"2863001c",
     8007 => x"f8000879",  8008 => x"78020001",  8009 => x"34010087",
     8010 => x"38424bd8",  8011 => x"f8000875",  8012 => x"29810000",
     8013 => x"b9601000",  8014 => x"28210020",  8015 => x"28240004",
     8016 => x"34010007",  8017 => x"28830028",  8018 => x"2884002c",
     8019 => x"f800086d",  8020 => x"e0000108",  8021 => x"78010001",
     8022 => x"38217594",  8023 => x"28210000",  8024 => x"34020001",
     8025 => x"4841000e",  8026 => x"34020002",  8027 => x"4c410004",
     8028 => x"34020003",  8029 => x"5c22000a",  8030 => x"e0000005",
     8031 => x"78020001",  8032 => x"34010007",  8033 => x"38424bf8",
     8034 => x"e0000008",  8035 => x"78020001",  8036 => x"34010007",
     8037 => x"38424c04",  8038 => x"e0000004",  8039 => x"78020001",
     8040 => x"34010001",  8041 => x"38424c10",  8042 => x"f8000856",
     8043 => x"2b810054",  8044 => x"44200005",  8045 => x"78020001",
     8046 => x"34010002",  8047 => x"38424c20",  8048 => x"e0000004",
     8049 => x"78020001",  8050 => x"34010001",  8051 => x"38424c2c",
     8052 => x"f800084c",  8053 => x"2b810070",  8054 => x"44200007",
     8055 => x"2b810074",  8056 => x"44200005",  8057 => x"78020001",
     8058 => x"34010002",  8059 => x"38424c38",  8060 => x"e0000004",
     8061 => x"78020001",  8062 => x"34010001",  8063 => x"38424c48",
     8064 => x"f8000840",  8065 => x"78020001",  8066 => x"38424c58",
     8067 => x"34010007",  8068 => x"f800083c",  8069 => x"378c0104",
     8070 => x"b9800800",  8071 => x"f8000bc8",  8072 => x"378300e8",
     8073 => x"b8600800",  8074 => x"b9801000",  8075 => x"5b83001c",
     8076 => x"f800069b",  8077 => x"78010001",  8078 => x"38217d90",
     8079 => x"28210000",  8080 => x"34020001",  8081 => x"2b83001c",
     8082 => x"4422000a",  8083 => x"44200004",  8084 => x"34020002",
     8085 => x"5c22000f",  8086 => x"e000000a",  8087 => x"78020001",
     8088 => x"34010001",  8089 => x"38424c60",  8090 => x"f8000826",
     8091 => x"e0000009",  8092 => x"78020001",  8093 => x"34010002",
     8094 => x"38424c70",  8095 => x"e0000004",  8096 => x"78020001",
     8097 => x"34010002",  8098 => x"38424c80",  8099 => x"f800081d",
     8100 => x"fbfffed9",  8101 => x"340d0001",  8102 => x"442000b6",
     8103 => x"78020001",  8104 => x"34010087",  8105 => x"38424c98",
     8106 => x"f8000816",  8107 => x"78020001",  8108 => x"34010007",
     8109 => x"38424860",  8110 => x"356300c0",  8111 => x"f8000811",
     8112 => x"78020001",  8113 => x"34010087",  8114 => x"38424cb4",
     8115 => x"f800080d",  8116 => x"296100bc",  8117 => x"44200005",
     8118 => x"78020001",  8119 => x"34010002",  8120 => x"38424cd0",
     8121 => x"e0000004",  8122 => x"78020001",  8123 => x"34010001",
     8124 => x"38424cd4",  8125 => x"f8000803",  8126 => x"78020001",
     8127 => x"34010087",  8128 => x"38424cdc",  8129 => x"f80007ff",
     8130 => x"34010000",  8131 => x"f800291e",  8132 => x"b8206000",
     8133 => x"20210001",  8134 => x"44200005",  8135 => x"78020001",
     8136 => x"34010002",  8137 => x"38424cf8",  8138 => x"f80007f6",
     8139 => x"218c0002",  8140 => x"45800005",  8141 => x"78020001",
     8142 => x"34010002",  8143 => x"38424d00",  8144 => x"f80007f0",
     8145 => x"78010001",  8146 => x"38214d20",  8147 => x"f800121c",
     8148 => x"78020001",  8149 => x"34010004",  8150 => x"38424d0c",
     8151 => x"f80007e9",  8152 => x"78020001",  8153 => x"34010087",
     8154 => x"38424d24",  8155 => x"f80007e5",  8156 => x"296200a4",
     8157 => x"296100a0",  8158 => x"780d0001",  8159 => x"39ad4d40",
     8160 => x"fbfffd9d",  8161 => x"b8201800",  8162 => x"b9a01000",
     8163 => x"34010007",  8164 => x"f80007dc",  8165 => x"78020001",
     8166 => x"34010087",  8167 => x"38424d48",  8168 => x"f80007d8",
     8169 => x"296200b4",  8170 => x"296100b0",  8171 => x"780c0001",
     8172 => x"398c4d80",  8173 => x"fbfffd90",  8174 => x"b8201800",
     8175 => x"b9a01000",  8176 => x"34010007",  8177 => x"f80007cf",
     8178 => x"78020001",  8179 => x"34010087",  8180 => x"38424d64",
     8181 => x"f80007cb",  8182 => x"29630018",  8183 => x"2964001c",
     8184 => x"b9801000",  8185 => x"34010007",  8186 => x"f80007c6",
     8187 => x"78020001",  8188 => x"34010087",  8189 => x"38424d98",
     8190 => x"f80007c2",  8191 => x"29640024",  8192 => x"29630020",
     8193 => x"b9801000",  8194 => x"34010007",  8195 => x"f80007bd",
     8196 => x"296e00b4",  8197 => x"296100a4",  8198 => x"78020001",
     8199 => x"3dce0001",  8200 => x"38424db4",  8201 => x"c82e7000",
     8202 => x"780c0001",  8203 => x"34010087",  8204 => x"f80007b4",
     8205 => x"398c4dd0",  8206 => x"b9c01800",  8207 => x"34010007",
     8208 => x"b9801000",  8209 => x"f80007af",  8210 => x"29610018",
     8211 => x"296200a4",  8212 => x"296f00a0",  8213 => x"1423001f",
     8214 => x"c8410800",  8215 => x"f4221000",  8216 => x"c9e37800",
     8217 => x"c9e27800",  8218 => x"2962001c",  8219 => x"296e0024",
     8220 => x"1443001f",  8221 => x"c8221000",  8222 => x"f4410800",
     8223 => x"c9e37800",  8224 => x"c9e17800",  8225 => x"29610020",
     8226 => x"1423001f",  8227 => x"c8410800",  8228 => x"f4221000",
     8229 => x"c9e37800",  8230 => x"15c3001f",  8231 => x"c82e7000",
     8232 => x"c9e27800",  8233 => x"f5c10800",  8234 => x"c9e37800",
     8235 => x"78020001",  8236 => x"c9e17800",  8237 => x"38424dd8",
     8238 => x"34010087",  8239 => x"f8000791",  8240 => x"b9c01000",
     8241 => x"b9e00800",  8242 => x"fbfffd4b",  8243 => x"b8201800",
     8244 => x"b9a01000",  8245 => x"34010007",  8246 => x"f800078a",
     8247 => x"78020001",  8248 => x"34010087",  8249 => x"38424df4",
     8250 => x"f8000786",  8251 => x"296300ec",  8252 => x"34010007",
     8253 => x"b9801000",  8254 => x"f8000782",  8255 => x"78020001",
     8256 => x"34010087",  8257 => x"38424e10",  8258 => x"f800077e",
     8259 => x"296300a8",  8260 => x"34010007",  8261 => x"b9801000",
     8262 => x"f800077a",  8263 => x"78020001",  8264 => x"34010087",
     8265 => x"38424e2c",  8266 => x"f8000776",  8267 => x"296300e4",
     8268 => x"34010007",  8269 => x"b9801000",  8270 => x"f8000772",
     8271 => x"78020001",  8272 => x"34010087",  8273 => x"38424e48",
     8274 => x"f800076e",  8275 => x"296300b8",  8276 => x"78020001",
     8277 => x"34010007",  8278 => x"38424e64",  8279 => x"f8000769",
     8280 => x"78010001",  8281 => x"38214e6c",  8282 => x"f8001195",
     8283 => x"340d0001",  8284 => x"b9a00800",  8285 => x"2b9d0004",
     8286 => x"2b8b0018",  8287 => x"2b8c0014",  8288 => x"2b8d0010",
     8289 => x"2b8e000c",  8290 => x"2b8f0008",  8291 => x"379c0110",
     8292 => x"c3a00000",  8293 => x"379cfff4",  8294 => x"5b8b0008",
     8295 => x"5b9d0004",  8296 => x"b8205800",  8297 => x"fbffe306",
     8298 => x"34020003",  8299 => x"5c220003",  8300 => x"34010002",
     8301 => x"e0000002",  8302 => x"34010001",  8303 => x"59610028",
     8304 => x"3562004c",  8305 => x"35610048",  8306 => x"f80012f8",
     8307 => x"34010000",  8308 => x"59600040",  8309 => x"59600044",
     8310 => x"59600088",  8311 => x"5960008c",  8312 => x"3782000c",
     8313 => x"34030000",  8314 => x"f80027dc",  8315 => x"44200006",
     8316 => x"2b81000c",  8317 => x"596100a0",  8318 => x"34010001",
     8319 => x"596100a4",  8320 => x"e0000003",  8321 => x"596000a0",
     8322 => x"596000a4",  8323 => x"34010000",  8324 => x"f80012be",
     8325 => x"5961002c",  8326 => x"34010001",  8327 => x"59610054",
     8328 => x"59610050",  8329 => x"34010000",  8330 => x"f8002767",
     8331 => x"59610034",  8332 => x"34011f40",  8333 => x"596100b4",
     8334 => x"78010001",  8335 => x"38216170",  8336 => x"28210000",
     8337 => x"596100b8",  8338 => x"596100bc",  8339 => x"35610014",
     8340 => x"f8001263",  8341 => x"34010000",  8342 => x"5960001c",
     8343 => x"2b9d0004",  8344 => x"2b8b0008",  8345 => x"379c000c",
     8346 => x"c3a00000",  8347 => x"c3a00000",  8348 => x"379cfffc",
     8349 => x"5b9d0004",  8350 => x"b8201000",  8351 => x"78010001",
     8352 => x"38214e80",  8353 => x"f800114e",  8354 => x"2b9d0004",
     8355 => x"379c0004",  8356 => x"c3a00000",  8357 => x"379cffcc",
     8358 => x"5b8b0010",  8359 => x"5b8c000c",  8360 => x"5b8d0008",
     8361 => x"5b9d0004",  8362 => x"378b0014",  8363 => x"34020000",
     8364 => x"34030024",  8365 => x"b9600800",  8366 => x"f8002b93",
     8367 => x"78030001",  8368 => x"b9600800",  8369 => x"34040000",
     8370 => x"34020000",  8371 => x"38637ac8",  8372 => x"34080020",
     8373 => x"34070008",  8374 => x"e0000004",  8375 => x"34840001",
     8376 => x"34210004",  8377 => x"44870017",  8378 => x"b4432800",
     8379 => x"e0000004",  8380 => x"30a00000",  8381 => x"34420001",
     8382 => x"34a50001",  8383 => x"40a60000",  8384 => x"44c8fffc",
     8385 => x"44c0000d",  8386 => x"b4432800",  8387 => x"58250000",
     8388 => x"e0000002",  8389 => x"34420001",  8390 => x"b4432800",
     8391 => x"40a50000",  8392 => x"7ca90000",  8393 => x"7ca60020",
     8394 => x"a1263000",  8395 => x"5cc0fffa",  8396 => x"5ca6ffeb",
     8397 => x"e0000003",  8398 => x"340c0000",  8399 => x"448c0021",
     8400 => x"2b810014",  8401 => x"340c0000",  8402 => x"40220000",
     8403 => x"34010023",  8404 => x"4441001c",  8405 => x"780b0001",
     8406 => x"780c0001",  8407 => x"396b7350",  8408 => x"398c7418",
     8409 => x"e0000011",  8410 => x"29610000",  8411 => x"f8002ba7",
     8412 => x"b8206800",  8413 => x"5c20000c",  8414 => x"29620004",
     8415 => x"37810018",  8416 => x"d8400000",  8417 => x"b8206000",
     8418 => x"4c2d000e",  8419 => x"29620000",  8420 => x"78010001",
     8421 => x"b9801800",  8422 => x"38214e88",  8423 => x"f8001108",
     8424 => x"e0000008",  8425 => x"356b0008",  8426 => x"2b820014",
     8427 => x"558bffef",  8428 => x"78010001",  8429 => x"38214ea0",
     8430 => x"f8001101",  8431 => x"340cffea",  8432 => x"b9800800",
     8433 => x"2b9d0004",  8434 => x"2b8b0010",  8435 => x"2b8c000c",
     8436 => x"2b8d0008",  8437 => x"379c0034",  8438 => x"c3a00000",
     8439 => x"379cfff8",  8440 => x"5b8b0008",  8441 => x"5b9d0004",
     8442 => x"780b0001",  8443 => x"396b7b1c",  8444 => x"29650000",
     8445 => x"78020001",  8446 => x"34240001",  8447 => x"b8201800",
     8448 => x"38427ac8",  8449 => x"b4220800",  8450 => x"c8a31800",
     8451 => x"b4821000",  8452 => x"f8002af8",  8453 => x"29610000",
     8454 => x"3421ffff",  8455 => x"59610000",  8456 => x"2b9d0004",
     8457 => x"2b8b0008",  8458 => x"379c0008",  8459 => x"c3a00000",
     8460 => x"78010001",  8461 => x"38217b24",  8462 => x"58200000",
     8463 => x"78010001",  8464 => x"38217b1c",  8465 => x"58200000",
     8466 => x"78010001",  8467 => x"38217b20",  8468 => x"58200000",
     8469 => x"c3a00000",  8470 => x"379cfff4",  8471 => x"5b8b000c",
     8472 => x"5b8c0008",  8473 => x"5b9d0004",  8474 => x"780b0001",
     8475 => x"396b7b20",  8476 => x"29610000",  8477 => x"340c0001",
     8478 => x"442c0010",  8479 => x"34020002",  8480 => x"4422009d",
     8481 => x"34020000",  8482 => x"5c2000a5",  8483 => x"78010001",
     8484 => x"38214ebc",  8485 => x"f80010ca",  8486 => x"78010001",
     8487 => x"38217b24",  8488 => x"58200000",  8489 => x"78010001",
     8490 => x"38217b1c",  8491 => x"58200000",  8492 => x"596c0000",
     8493 => x"e000008e",  8494 => x"f8002104",  8495 => x"34020000",
     8496 => x"48010097",  8497 => x"3402001b",  8498 => x"44220008",
     8499 => x"78020001",  8500 => x"38427b28",  8501 => x"28430000",
     8502 => x"6424005b",  8503 => x"00650010",  8504 => x"a0a42000",
     8505 => x"44800006",  8506 => x"78010001",  8507 => x"38217b28",
     8508 => x"78020001",  8509 => x"58220000",  8510 => x"e0000003",
     8511 => x"b8230800",  8512 => x"58410000",  8513 => x"78010001",
     8514 => x"38217b28",  8515 => x"282b0000",  8516 => x"34020001",
     8517 => x"216100ff",  8518 => x"44200081",  8519 => x"3401007e",
     8520 => x"4561002e",  8521 => x"49610006",  8522 => x"34010009",
     8523 => x"4561006d",  8524 => x"3401000d",  8525 => x"5d610042",
     8526 => x"e0000020",  8527 => x"78020001",  8528 => x"38425a58",
     8529 => x"28410000",  8530 => x"45610010",  8531 => x"78020001",
     8532 => x"38425a5c",  8533 => x"28410000",  8534 => x"45610004",
     8535 => x"3401007f",  8536 => x"5d610037",  8537 => x"e0000027",
     8538 => x"78010001",  8539 => x"38217b24",  8540 => x"28220000",
     8541 => x"4c02005b",  8542 => x"3442ffff",  8543 => x"58220000",
     8544 => x"34010044",  8545 => x"e000000b",  8546 => x"78010001",
     8547 => x"78020001",  8548 => x"38217b24",  8549 => x"38427b1c",
     8550 => x"28230000",  8551 => x"28420000",  8552 => x"4c620050",
     8553 => x"34630001",  8554 => x"58230000",  8555 => x"34010043",
     8556 => x"fbffff30",  8557 => x"e000004b",  8558 => x"78010001",
     8559 => x"38214d20",  8560 => x"f800107f",  8561 => x"78010001",
     8562 => x"38217b20",  8563 => x"34020002",  8564 => x"58220000",
     8565 => x"e0000043",  8566 => x"78010001",  8567 => x"78020001",
     8568 => x"38217b24",  8569 => x"38427b1c",  8570 => x"28210000",
     8571 => x"28420000",  8572 => x"4422003c",  8573 => x"fbffff7a",
     8574 => x"34010050",  8575 => x"e3ffffed",  8576 => x"780b0001",
     8577 => x"396b7b24",  8578 => x"29610000",  8579 => x"4c010035",
     8580 => x"34010044",  8581 => x"fbffff17",  8582 => x"34010050",
     8583 => x"fbffff15",  8584 => x"29610000",  8585 => x"3421ffff",
     8586 => x"fbffff6d",  8587 => x"29610000",  8588 => x"3421ffff",
     8589 => x"59610000",  8590 => x"e000002a",  8591 => x"78010001",
     8592 => x"a1610800",  8593 => x"5c200027",  8594 => x"78010001",
     8595 => x"38217b1c",  8596 => x"28240000",  8597 => x"3401004f",
     8598 => x"48810022",  8599 => x"78010001",  8600 => x"38217b24",
     8601 => x"28230000",  8602 => x"44640008",  8603 => x"78020001",
     8604 => x"34610001",  8605 => x"38427ac8",  8606 => x"b4220800",
     8607 => x"b4621000",  8608 => x"c8831800",  8609 => x"f8002a5b",
     8610 => x"78010001",  8611 => x"38217b24",  8612 => x"28230000",
     8613 => x"78020001",  8614 => x"38427ac8",  8615 => x"b4431000",
     8616 => x"304b0000",  8617 => x"34620001",  8618 => x"58220000",
     8619 => x"78010001",  8620 => x"38217b1c",  8621 => x"28220000",
     8622 => x"34420001",  8623 => x"58220000",  8624 => x"34010040",
     8625 => x"fbfffeeb",  8626 => x"78020001",  8627 => x"38427b28",
     8628 => x"28420000",  8629 => x"78010001",  8630 => x"38214ec4",
     8631 => x"f8001038",  8632 => x"78010001",  8633 => x"38217b28",
     8634 => x"58200000",  8635 => x"34020001",  8636 => x"e000000b",
     8637 => x"78020001",  8638 => x"38427b1c",  8639 => x"28420000",
     8640 => x"78010001",  8641 => x"38217ac8",  8642 => x"b4220800",
     8643 => x"30200000",  8644 => x"fbfffee1",  8645 => x"59600000",
     8646 => x"e3fffff5",  8647 => x"b8400800",  8648 => x"2b9d0004",
     8649 => x"2b8b000c",  8650 => x"2b8c0008",  8651 => x"379c000c",
     8652 => x"c3a00000",  8653 => x"34030000",  8654 => x"34070009",
     8655 => x"34050005",  8656 => x"e0000014",  8657 => x"3486ffd0",
     8658 => x"20c800ff",  8659 => x"55070004",  8660 => x"3c630004",
     8661 => x"b4c31800",  8662 => x"e000000d",  8663 => x"3486ffbf",
     8664 => x"20c600ff",  8665 => x"54c50004",  8666 => x"3c630004",
     8667 => x"3484ffc9",  8668 => x"e0000006",  8669 => x"3486ff9f",
     8670 => x"20c600ff",  8671 => x"54c50007",  8672 => x"3c630004",
     8673 => x"3484ffa9",  8674 => x"b4831800",  8675 => x"34210001",
     8676 => x"40240000",  8677 => x"5c80ffec",  8678 => x"58430000",
     8679 => x"c3a00000",  8680 => x"34030000",  8681 => x"34050009",
     8682 => x"e0000007",  8683 => x"3484ffd0",  8684 => x"208600ff",
     8685 => x"54c50006",  8686 => x"0863000a",  8687 => x"34210001",
     8688 => x"b4831800",  8689 => x"40240000",  8690 => x"5c80fff9",
     8691 => x"58430000",  8692 => x"c3a00000",  8693 => x"379cffec",
     8694 => x"5b8b0014",  8695 => x"5b8c0010",  8696 => x"5b8d000c",
     8697 => x"5b8e0008",  8698 => x"5b9d0004",  8699 => x"78010001",
     8700 => x"38218efc",  8701 => x"40210000",  8702 => x"4420001b",
     8703 => x"780b0001",  8704 => x"780e0001",  8705 => x"780d0001",
     8706 => x"340c0000",  8707 => x"396b7ac8",  8708 => x"39ce7b1c",
     8709 => x"39ad4ee0",  8710 => x"b9600800",  8711 => x"34020050",
     8712 => x"b9801800",  8713 => x"f8001c1a",  8714 => x"59c10000",
     8715 => x"48200006",  8716 => x"5d80000d",  8717 => x"78010001",
     8718 => x"38214ec8",  8719 => x"f8000fe0",  8720 => x"e0000009",
     8721 => x"b5610800",  8722 => x"3020ffff",  8723 => x"b9601000",
     8724 => x"b9a00800",  8725 => x"f8000fda",  8726 => x"fbfffe8f",
     8727 => x"340c0001",  8728 => x"e3ffffee",  8729 => x"2b9d0004",
     8730 => x"2b8b0014",  8731 => x"2b8c0010",  8732 => x"2b8d000c",
     8733 => x"2b8e0008",  8734 => x"379c0014",  8735 => x"c3a00000",
     8736 => x"379cfff8",  8737 => x"5b8b0008",  8738 => x"5b9d0004",
     8739 => x"78010001",  8740 => x"382192a8",  8741 => x"28210000",
     8742 => x"78030001",  8743 => x"38636158",  8744 => x"28620000",
     8745 => x"282b000c",  8746 => x"78030001",  8747 => x"78010001",
     8748 => x"38634f08",  8749 => x"38214ef0",  8750 => x"f8000fc1",
     8751 => x"78050001",  8752 => x"78030001",  8753 => x"78040001",
     8754 => x"38a5615c",  8755 => x"38636160",  8756 => x"38846164",
     8757 => x"28a20000",  8758 => x"28630000",  8759 => x"28840000",
     8760 => x"78010001",  8761 => x"38214f28",  8762 => x"f8000fb5",
     8763 => x"216b000f",  8764 => x"356b0001",  8765 => x"78010001",
     8766 => x"34020080",  8767 => x"3d6b0004",  8768 => x"38214f3c",
     8769 => x"34030800",  8770 => x"f8000fad",  8771 => x"3561ff80",
     8772 => x"3402000f",  8773 => x"50410006",  8774 => x"78010001",
     8775 => x"38214f64",  8776 => x"b9601000",  8777 => x"35630010",
     8778 => x"f8000fa5",  8779 => x"34010000",  8780 => x"2b9d0004",
     8781 => x"2b8b0008",  8782 => x"379c0008",  8783 => x"c3a00000",
     8784 => x"379cfff8",  8785 => x"5b8b0008",  8786 => x"5b9d0004",
     8787 => x"b8205800",  8788 => x"28210000",  8789 => x"78020001",
     8790 => x"38424f94",  8791 => x"f8002a2b",  8792 => x"5c200003",
     8793 => x"fbffe11a",  8794 => x"e0000008",  8795 => x"29610000",
     8796 => x"78020001",  8797 => x"38424f9c",  8798 => x"f8002a24",
     8799 => x"3402ffea",  8800 => x"5c200003",  8801 => x"fbffe138",
     8802 => x"b8201000",  8803 => x"b8400800",  8804 => x"2b9d0004",
     8805 => x"2b8b0008",  8806 => x"379c0008",  8807 => x"c3a00000",
     8808 => x"379cfff8",  8809 => x"5b8b0008",  8810 => x"5b9d0004",
     8811 => x"b8205800",  8812 => x"28210000",  8813 => x"78020001",
     8814 => x"38424fa4",  8815 => x"f8002a13",  8816 => x"34020001",
     8817 => x"44200018",  8818 => x"29610000",  8819 => x"78020001",
     8820 => x"3842435c",  8821 => x"f8002a0d",  8822 => x"34020002",
     8823 => x"44200012",  8824 => x"29610000",  8825 => x"78020001",
     8826 => x"38423e74",  8827 => x"f8002a07",  8828 => x"34020003",
     8829 => x"4420000c",  8830 => x"fbffe0f1",  8831 => x"3c210002",
     8832 => x"78020001",  8833 => x"38425d38",  8834 => x"b4411000",
     8835 => x"28420000",  8836 => x"78010001",  8837 => x"38214860",
     8838 => x"f8000f69",  8839 => x"34010000",  8840 => x"e0000003",
     8841 => x"b8400800",  8842 => x"fbffe135",  8843 => x"2b9d0004",
     8844 => x"2b8b0008",  8845 => x"379c0008",  8846 => x"c3a00000",
     8847 => x"379cfff0",  8848 => x"5b8b0010",  8849 => x"5b8c000c",
     8850 => x"5b8d0008",  8851 => x"5b9d0004",  8852 => x"78010001",
     8853 => x"38214fbc",  8854 => x"780b0001",  8855 => x"780d0001",
     8856 => x"780c0001",  8857 => x"f8000f56",  8858 => x"396b7350",
     8859 => x"39ad7418",  8860 => x"398c4fd4",  8861 => x"e0000005",
     8862 => x"29620000",  8863 => x"b9800800",  8864 => x"356b0008",
     8865 => x"f8000f4e",  8866 => x"55abfffc",  8867 => x"34010000",
     8868 => x"2b9d0004",  8869 => x"2b8b0010",  8870 => x"2b8c000c",
     8871 => x"2b8d0008",  8872 => x"379c0010",  8873 => x"c3a00000",
     8874 => x"379cffec",  8875 => x"5b8b0010",  8876 => x"5b8c000c",
     8877 => x"5b8d0008",  8878 => x"5b9d0004",  8879 => x"340b0000",
     8880 => x"b8406800",  8881 => x"340c0006",  8882 => x"37820014",
     8883 => x"fbffff1a",  8884 => x"2b830014",  8885 => x"b5ab1000",
     8886 => x"356b0001",  8887 => x"30430000",  8888 => x"40220000",
     8889 => x"6442003a",  8890 => x"b4220800",  8891 => x"5d6cfff7",
     8892 => x"2b9d0004",  8893 => x"2b8b0010",  8894 => x"2b8c000c",
     8895 => x"2b8d0008",  8896 => x"379c0014",  8897 => x"c3a00000",
     8898 => x"379cfff8",  8899 => x"5b8b0008",  8900 => x"5b9d0004",
     8901 => x"b8404000",  8902 => x"41030000",  8903 => x"41040001",
     8904 => x"41050002",  8905 => x"41060003",  8906 => x"41070004",
     8907 => x"41080005",  8908 => x"78020001",  8909 => x"38424fe4",
     8910 => x"b8205800",  8911 => x"f8000f12",  8912 => x"b9600800",
     8913 => x"2b9d0004",  8914 => x"2b8b0008",  8915 => x"379c0008",
     8916 => x"c3a00000",  8917 => x"379cffd0",  8918 => x"5b8b0008",
     8919 => x"5b9d0004",  8920 => x"b8205800",  8921 => x"28210000",
     8922 => x"44200005",  8923 => x"78020001",  8924 => x"38425004",
     8925 => x"f80029a5",  8926 => x"5c200004",  8927 => x"3781002c",
     8928 => x"f8001017",  8929 => x"e000002b",  8930 => x"29610000",
     8931 => x"78020001",  8932 => x"38425008",  8933 => x"f800299d",
     8934 => x"5c200008",  8935 => x"378b002c",  8936 => x"b9600800",
     8937 => x"f800100e",  8938 => x"b9601000",  8939 => x"34010000",
     8940 => x"f8001b92",  8941 => x"e000001f",  8942 => x"29610000",
     8943 => x"78020001",  8944 => x"38425010",  8945 => x"f8002991",
     8946 => x"5c20000b",  8947 => x"29630004",  8948 => x"44610009",
     8949 => x"378b002c",  8950 => x"b8600800",  8951 => x"b9601000",
     8952 => x"fbffffb2",  8953 => x"b9600800",  8954 => x"f8000fe9",
     8955 => x"f80010e4",  8956 => x"e0000010",  8957 => x"29610000",
     8958 => x"78020001",  8959 => x"38425014",  8960 => x"f8002982",
     8961 => x"b8201800",  8962 => x"3402ffea",  8963 => x"5c200011",
     8964 => x"29610004",  8965 => x"4423000f",  8966 => x"378b002c",
     8967 => x"b9601000",  8968 => x"fbffffa2",  8969 => x"34010000",
     8970 => x"b9601000",  8971 => x"f8001b6a",  8972 => x"3782002c",
     8973 => x"3781000c",  8974 => x"fbffffb4",  8975 => x"b8201000",
     8976 => x"78010001",  8977 => x"3821501c",  8978 => x"f8000edd",
     8979 => x"34020000",  8980 => x"b8400800",  8981 => x"2b9d0004",
     8982 => x"2b8b0008",  8983 => x"379c0030",  8984 => x"c3a00000",
     8985 => x"379cffe8",  8986 => x"5b8b0018",  8987 => x"5b8c0014",
     8988 => x"5b8d0010",  8989 => x"5b8e000c",  8990 => x"5b8f0008",
     8991 => x"5b9d0004",  8992 => x"28210000",  8993 => x"44200010",
     8994 => x"78020001",  8995 => x"38425034",  8996 => x"f800295e",
     8997 => x"5c20000c",  8998 => x"78010001",  8999 => x"78020001",
     9000 => x"38217424",  9001 => x"38427574",  9002 => x"e0000005",
     9003 => x"58200018",  9004 => x"58200014",  9005 => x"58200010",
     9006 => x"3421001c",  9007 => x"5441fffc",  9008 => x"e0000018",
     9009 => x"78010001",  9010 => x"3821503c",  9011 => x"780b0001",
     9012 => x"780d0001",  9013 => x"780c0001",  9014 => x"f8000eb9",
     9015 => x"396b7424",  9016 => x"39ad7574",  9017 => x"398c5064",
     9018 => x"e000000d",  9019 => x"29610018",  9020 => x"340203e8",
     9021 => x"296f0010",  9022 => x"f8002824",  9023 => x"296e0014",
     9024 => x"29650000",  9025 => x"b8202000",  9026 => x"b9e01000",
     9027 => x"b9800800",  9028 => x"b9c01800",  9029 => x"f8000eaa",
     9030 => x"356b001c",  9031 => x"55abfff4",  9032 => x"34010000",
     9033 => x"2b9d0004",  9034 => x"2b8b0018",  9035 => x"2b8c0014",
     9036 => x"2b8d0010",  9037 => x"2b8e000c",  9038 => x"2b8f0008",
     9039 => x"379c0018",  9040 => x"c3a00000",  9041 => x"379cfff8",
     9042 => x"5b9d0004",  9043 => x"b8201000",  9044 => x"28210000",
     9045 => x"4420000d",  9046 => x"28420004",  9047 => x"5c40000b",
     9048 => x"37820008",  9049 => x"fbfffe8f",  9050 => x"2b820008",
     9051 => x"78010001",  9052 => x"38216168",  9053 => x"084203e8",
     9054 => x"58220000",  9055 => x"78010001",  9056 => x"38214d20",
     9057 => x"e0000003",  9058 => x"78010001",  9059 => x"38215084",
     9060 => x"f8000e8b",  9061 => x"34010000",  9062 => x"2b9d0004",
     9063 => x"379c0008",  9064 => x"c3a00000",  9065 => x"379cfff8",
     9066 => x"5b8b0008",  9067 => x"5b9d0004",  9068 => x"b8205800",
     9069 => x"28210000",  9070 => x"5c200011",  9071 => x"78010001",
     9072 => x"38219290",  9073 => x"28220000",  9074 => x"340b0000",
     9075 => x"64420000",  9076 => x"58220000",  9077 => x"78010001",
     9078 => x"38218f2c",  9079 => x"28230000",  9080 => x"3463ffff",
     9081 => x"58230000",  9082 => x"5c4b002b",  9083 => x"78010001",
     9084 => x"382150a8",  9085 => x"f8000e72",  9086 => x"e0000027",
     9087 => x"78020001",  9088 => x"384250bc",  9089 => x"f8002901",
     9090 => x"5c200007",  9091 => x"f8000fdd",  9092 => x"b8201000",
     9093 => x"78010001",  9094 => x"38215790",  9095 => x"f8000e68",
     9096 => x"e000001c",  9097 => x"29610000",  9098 => x"78020001",
     9099 => x"38423f14",  9100 => x"f80028f6",  9101 => x"5c20000b",
     9102 => x"78010001",  9103 => x"38219290",  9104 => x"34020001",
     9105 => x"58220000",  9106 => x"78010001",  9107 => x"38218f2c",
     9108 => x"28220000",  9109 => x"3442ffff",  9110 => x"58220000",
     9111 => x"e000000d",  9112 => x"29610000",  9113 => x"78020001",
     9114 => x"384250c0",  9115 => x"f80028e7",  9116 => x"340bffea",
     9117 => x"5c200008",  9118 => x"78010001",  9119 => x"38219290",
     9120 => x"58200000",  9121 => x"78010001",  9122 => x"382150a8",
     9123 => x"f8000e4c",  9124 => x"340b0000",  9125 => x"b9600800",
     9126 => x"2b9d0004",  9127 => x"2b8b0008",  9128 => x"379c0008",
     9129 => x"c3a00000",  9130 => x"379cffb8",  9131 => x"5b8b0028",
     9132 => x"5b8c0024",  9133 => x"5b8d0020",  9134 => x"5b8e001c",
     9135 => x"5b8f0018",  9136 => x"5b900014",  9137 => x"5b910010",
     9138 => x"5b92000c",  9139 => x"5b930008",  9140 => x"5b9d0004",
     9141 => x"b8205800",  9142 => x"28210000",  9143 => x"442000c8",
     9144 => x"78020001",  9145 => x"384250e0",  9146 => x"f80028c8",
     9147 => x"5c200008",  9148 => x"f8001870",  9149 => x"3403ffff",
     9150 => x"34020000",  9151 => x"5c2300c4",  9152 => x"78010001",
     9153 => x"382150e8",  9154 => x"e000003c",  9155 => x"29610010",
     9156 => x"44200045",  9157 => x"29610000",  9158 => x"78020001",
     9159 => x"384250fc",  9160 => x"f80028ba",  9161 => x"5c200040",
     9162 => x"29610004",  9163 => x"34020010",  9164 => x"356c0004",
     9165 => x"f80029d9",  9166 => x"3c210018",  9167 => x"34030000",
     9168 => x"14210018",  9169 => x"3784002c",  9170 => x"e0000007",
     9171 => x"29820000",  9172 => x"b4832800",  9173 => x"b4431000",
     9174 => x"40420000",  9175 => x"34630001",  9176 => x"30a20000",
     9177 => x"b0601000",  9178 => x"4822fff9",  9179 => x"b4820800",
     9180 => x"34030020",  9181 => x"3404000f",  9182 => x"e0000005",
     9183 => x"34420001",  9184 => x"30230000",  9185 => x"b0401000",
     9186 => x"34210001",  9187 => x"4c82fffc",  9188 => x"29610008",
     9189 => x"f8000429",  9190 => x"5b810040",  9191 => x"2961000c",
     9192 => x"f8000426",  9193 => x"5b810044",  9194 => x"29610010",
     9195 => x"f8000423",  9196 => x"5b81003c",  9197 => x"34020001",
     9198 => x"3781002c",  9199 => x"34030000",  9200 => x"f8001855",
     9201 => x"3c220018",  9202 => x"3401fffe",  9203 => x"14420018",
     9204 => x"5c410006",  9205 => x"78010001",  9206 => x"38215100",
     9207 => x"f8000df8",  9208 => x"3402ffe4",  9209 => x"e000008a",
     9210 => x"3401ffff",  9211 => x"5c410006",  9212 => x"78010001",
     9213 => x"38215110",  9214 => x"f8000df1",  9215 => x"3402fffb",
     9216 => x"e0000083",  9217 => x"4c400004",  9218 => x"78010001",
     9219 => x"3821511c",  9220 => x"e0000023",  9221 => x"78010001",
     9222 => x"38215138",  9223 => x"f8000de8",  9224 => x"e0000075",
     9225 => x"29610000",  9226 => x"78020001",  9227 => x"38425148",
     9228 => x"f8002876",  9229 => x"5c200030",  9230 => x"78100001",
     9231 => x"780f0001",  9232 => x"780e0001",  9233 => x"340c0000",
     9234 => x"34110000",  9235 => x"3792002c",  9236 => x"3a105164",
     9237 => x"3793003c",  9238 => x"39ef4ec4",  9239 => x"39ce516c",
     9240 => x"ba400800",  9241 => x"34020000",  9242 => x"b9801800",
     9243 => x"f800182a",  9244 => x"3c2b0018",  9245 => x"156b0018",
     9246 => x"5d600005",  9247 => x"78010001",  9248 => x"38215150",
     9249 => x"f8000dce",  9250 => x"e000005b",  9251 => x"4d600007",
     9252 => x"78010001",  9253 => x"3821511c",  9254 => x"b9601000",
     9255 => x"f8000dc8",  9256 => x"3402fff2",  9257 => x"e000005a",
     9258 => x"358c0001",  9259 => x"ba000800",  9260 => x"b9801000",
     9261 => x"f8000dc2",  9262 => x"ba406800",  9263 => x"41a20000",
     9264 => x"b9e00800",  9265 => x"35ad0001",  9266 => x"f8000dbd",
     9267 => x"5db3fffc",  9268 => x"2b820040",  9269 => x"2b830044",
     9270 => x"2b84003c",  9271 => x"36310001",  9272 => x"b9c00800",
     9273 => x"b2208800",  9274 => x"f8000db5",  9275 => x"4971ffdd",
     9276 => x"e0000041",  9277 => x"29610000",  9278 => x"78020001",
     9279 => x"3842518c",  9280 => x"f8002842",  9281 => x"5c200032",
     9282 => x"f80013c8",  9283 => x"3c2c0018",  9284 => x"3401ffed",
     9285 => x"158c0018",  9286 => x"5d810006",  9287 => x"78010001",
     9288 => x"38215194",  9289 => x"f8000da6",  9290 => x"3402ffed",
     9291 => x"e0000038",  9292 => x"780b0001",  9293 => x"396b8f34",
     9294 => x"780d0001",  9295 => x"3401fffb",  9296 => x"356e0010",
     9297 => x"39ad4ec4",  9298 => x"5d810004",  9299 => x"78010001",
     9300 => x"382151a0",  9301 => x"e3ffffa9",  9302 => x"41620000",
     9303 => x"b9a00800",  9304 => x"356b0001",  9305 => x"f8000d96",
     9306 => x"5d6efffc",  9307 => x"78010001",  9308 => x"38214d20",
     9309 => x"f8000d92",  9310 => x"3401fffa",  9311 => x"5d810006",
     9312 => x"78010001",  9313 => x"382151b0",  9314 => x"f8000d8d",
     9315 => x"3402fffa",  9316 => x"e000001f",  9317 => x"78020001",
     9318 => x"78030001",  9319 => x"78040001",  9320 => x"38428ec8",
     9321 => x"38638ecc",  9322 => x"38846ffc",  9323 => x"28420000",
     9324 => x"28630000",  9325 => x"28840000",  9326 => x"78010001",
     9327 => x"382151c8",  9328 => x"f8000d7f",  9329 => x"b9801000",
     9330 => x"e0000011",  9331 => x"29610004",  9332 => x"4420000b",
     9333 => x"29610000",  9334 => x"78020001",  9335 => x"384251f0",
     9336 => x"f800280a",  9337 => x"5c200006",  9338 => x"29610004",
     9339 => x"f8000393",  9340 => x"f8000f31",  9341 => x"34020000",
     9342 => x"e0000005",  9343 => x"78010001",  9344 => x"382150cc",
     9345 => x"f8000d6e",  9346 => x"3402ffea",  9347 => x"b8400800",
     9348 => x"2b9d0004",  9349 => x"2b8b0028",  9350 => x"2b8c0024",
     9351 => x"2b8d0020",  9352 => x"2b8e001c",  9353 => x"2b8f0018",
     9354 => x"2b900014",  9355 => x"2b910010",  9356 => x"2b92000c",
     9357 => x"2b930008",  9358 => x"379c0048",  9359 => x"c3a00000",
     9360 => x"379cffe8",  9361 => x"5b8b0010",  9362 => x"5b8c000c",
     9363 => x"5b8d0008",  9364 => x"5b9d0004",  9365 => x"b8205800",
     9366 => x"28210000",  9367 => x"78020001",  9368 => x"384251f8",
     9369 => x"f80027e9",  9370 => x"5c200011",  9371 => x"2963000c",
     9372 => x"3402ffea",  9373 => x"44610086",  9374 => x"29610004",
     9375 => x"f800036f",  9376 => x"b8206800",  9377 => x"29610008",
     9378 => x"f800036c",  9379 => x"b8206000",  9380 => x"2961000c",
     9381 => x"f8000369",  9382 => x"b8201800",  9383 => x"b9801000",
     9384 => x"b9a00800",  9385 => x"f800227e",  9386 => x"e0000078",
     9387 => x"29610000",  9388 => x"78020001",  9389 => x"38425200",
     9390 => x"f80027d4",  9391 => x"b8201800",  9392 => x"5c200007",
     9393 => x"29610004",  9394 => x"3402ffea",  9395 => x"44230070",
     9396 => x"f800035a",  9397 => x"f800233c",  9398 => x"e0000060",
     9399 => x"29610000",  9400 => x"78020001",  9401 => x"384250c4",
     9402 => x"f80027c8",  9403 => x"5c200003",  9404 => x"f80023cf",
     9405 => x"e0000065",  9406 => x"29610000",  9407 => x"78020001",
     9408 => x"38425204",  9409 => x"f80027c1",  9410 => x"5c20000d",
     9411 => x"29630008",  9412 => x"3402ffea",  9413 => x"4461005e",
     9414 => x"29610004",  9415 => x"f8000347",  9416 => x"b8206000",
     9417 => x"29610008",  9418 => x"f8000344",  9419 => x"b8201000",
     9420 => x"b9800800",  9421 => x"f8002335",  9422 => x"e0000054",
     9423 => x"29610000",  9424 => x"78020001",  9425 => x"38425208",
     9426 => x"f80027b0",  9427 => x"b8201800",  9428 => x"5c20000e",
     9429 => x"29610004",  9430 => x"3402ffea",  9431 => x"4423004c",
     9432 => x"f8000336",  9433 => x"37820018",  9434 => x"37830014",
     9435 => x"f800234f",  9436 => x"2b820018",  9437 => x"2b830014",
     9438 => x"78010001",  9439 => x"3821520c",  9440 => x"f8000d0f",
     9441 => x"e0000041",  9442 => x"29610000",  9443 => x"78020001",
     9444 => x"38424f94",  9445 => x"f800279d",  9446 => x"b8201800",
     9447 => x"5c200007",  9448 => x"29610004",  9449 => x"3402ffea",
     9450 => x"44230039",  9451 => x"f8000323",  9452 => x"f80022e7",
     9453 => x"e0000035",  9454 => x"29610000",  9455 => x"78020001",
     9456 => x"38424f9c",  9457 => x"f8002791",  9458 => x"b8201800",
     9459 => x"5c200007",  9460 => x"29610004",  9461 => x"3402ffea",
     9462 => x"4423002d",  9463 => x"f8000317",  9464 => x"f80022ec",
     9465 => x"e0000029",  9466 => x"29610000",  9467 => x"78020001",
     9468 => x"38425214",  9469 => x"f8002785",  9470 => x"5c20000d",
     9471 => x"29630008",  9472 => x"3402ffea",  9473 => x"44610022",
     9474 => x"29610004",  9475 => x"f800030b",  9476 => x"b8206000",
     9477 => x"29610008",  9478 => x"f8000308",  9479 => x"b8201000",
     9480 => x"b9800800",  9481 => x"f80023f2",  9482 => x"e0000018",
     9483 => x"29610000",  9484 => x"78020001",  9485 => x"3842521c",
     9486 => x"f8002774",  9487 => x"b8201800",  9488 => x"5c20000b",
     9489 => x"29610004",  9490 => x"3402ffea",  9491 => x"44230010",
     9492 => x"f80002fa",  9493 => x"f80023d7",  9494 => x"b8201000",
     9495 => x"78010001",  9496 => x"38214e9c",  9497 => x"f8000cd6",
     9498 => x"e0000008",  9499 => x"29610000",  9500 => x"78020001",
     9501 => x"38425224",  9502 => x"f8002764",  9503 => x"3402ffea",
     9504 => x"5c200003",  9505 => x"f8002489",  9506 => x"34020000",
     9507 => x"b8400800",  9508 => x"2b9d0004",  9509 => x"2b8b0010",
     9510 => x"2b8c000c",  9511 => x"2b8d0008",  9512 => x"379c0018",
     9513 => x"c3a00000",  9514 => x"379cfff0",  9515 => x"5b8b000c",
     9516 => x"5b8c0008",  9517 => x"5b9d0004",  9518 => x"b8205800",
     9519 => x"28210000",  9520 => x"4420000b",  9521 => x"78020001",
     9522 => x"38425234",  9523 => x"f800274f",  9524 => x"b8206000",
     9525 => x"5c200006",  9526 => x"37810010",  9527 => x"f800141e",
     9528 => x"340bffff",  9529 => x"49810021",  9530 => x"e000001c",
     9531 => x"29610000",  9532 => x"340b0000",  9533 => x"5c20001d",
     9534 => x"37810010",  9535 => x"34020000",  9536 => x"f80017de",
     9537 => x"4d61000a",  9538 => x"2b820010",  9539 => x"78010001",
     9540 => x"3821523c",  9541 => x"f8000caa",  9542 => x"2b820010",
     9543 => x"78010001",  9544 => x"38216170",  9545 => x"58220000",
     9546 => x"e0000010",  9547 => x"78010001",  9548 => x"38215264",
     9549 => x"f8000ca2",  9550 => x"37810010",  9551 => x"f8001406",
     9552 => x"340bffff",  9553 => x"48010009",  9554 => x"2b820010",
     9555 => x"78010001",  9556 => x"38216170",  9557 => x"58220000",
     9558 => x"37810010",  9559 => x"34020001",  9560 => x"f80017c6",
     9561 => x"b8205800",  9562 => x"b9600800",  9563 => x"2b9d0004",
     9564 => x"2b8b000c",  9565 => x"2b8c0008",  9566 => x"379c0010",
     9567 => x"c3a00000",  9568 => x"379cffe8",  9569 => x"5b8b000c",
     9570 => x"5b8c0008",  9571 => x"5b9d0004",  9572 => x"b8205800",
     9573 => x"37820018",  9574 => x"37810010",  9575 => x"f80015e4",
     9576 => x"29610008",  9577 => x"44200014",  9578 => x"29610000",
     9579 => x"78020001",  9580 => x"38425010",  9581 => x"f8002715",
     9582 => x"5c20000f",  9583 => x"fbffde00",  9584 => x"34030003",
     9585 => x"3402fff0",  9586 => x"44230040",  9587 => x"29610004",
     9588 => x"f800029a",  9589 => x"b8206000",  9590 => x"29610008",
     9591 => x"f8000297",  9592 => x"b8201800",  9593 => x"b9801000",
     9594 => x"1581001f",  9595 => x"34040003",  9596 => x"e0000020",
     9597 => x"29610000",  9598 => x"4420000f",  9599 => x"78020001",
     9600 => x"38425298",  9601 => x"f8002701",  9602 => x"5c20000b",
     9603 => x"fbffddec",  9604 => x"34020003",  9605 => x"44220023",
     9606 => x"29610004",  9607 => x"f8000287",  9608 => x"b8201000",
     9609 => x"34030000",  9610 => x"1421001f",  9611 => x"34040001",
     9612 => x"e0000010",  9613 => x"29610000",  9614 => x"44200010",
     9615 => x"78020001",  9616 => x"384252a0",  9617 => x"f80026f1",
     9618 => x"5c20000c",  9619 => x"fbffdddc",  9620 => x"34020003",
     9621 => x"44220013",  9622 => x"29610004",  9623 => x"f8000277",
     9624 => x"b8201800",  9625 => x"34020000",  9626 => x"34010000",
     9627 => x"34040002",  9628 => x"f800158f",  9629 => x"e0000014",
     9630 => x"29610000",  9631 => x"44200009",  9632 => x"78020001",
     9633 => x"384252a8",  9634 => x"f80026e0",  9635 => x"5c200005",
     9636 => x"78010001",  9637 => x"3821520c",  9638 => x"2b820014",
     9639 => x"e0000008",  9640 => x"2b820014",  9641 => x"2b810010",
     9642 => x"34030000",  9643 => x"f8000164",  9644 => x"b8201000",
     9645 => x"78010001",  9646 => x"382152ac",  9647 => x"2b830018",
     9648 => x"f8000c3f",  9649 => x"34020000",  9650 => x"b8400800",
     9651 => x"2b9d0004",  9652 => x"2b8b000c",  9653 => x"2b8c0008",
     9654 => x"379c0018",  9655 => x"c3a00000",  9656 => x"78010001",
     9657 => x"38217578",  9658 => x"34020001",  9659 => x"58220000",
     9660 => x"34010000",  9661 => x"c3a00000",  9662 => x"379cfffc",
     9663 => x"5b9d0004",  9664 => x"f800127e",  9665 => x"34010000",
     9666 => x"2b9d0004",  9667 => x"379c0004",  9668 => x"c3a00000",
     9669 => x"379cfff8",  9670 => x"5b8b0008",  9671 => x"5b9d0004",
     9672 => x"b8205800",  9673 => x"28210000",  9674 => x"4420000c",
     9675 => x"78020001",  9676 => x"384252dc",  9677 => x"f80026b5",
     9678 => x"5c200008",  9679 => x"34010001",  9680 => x"fbffe890",
     9681 => x"78010001",  9682 => x"3821616c",  9683 => x"34020001",
     9684 => x"58220000",  9685 => x"e000000b",  9686 => x"29610000",
     9687 => x"44200009",  9688 => x"78020001",  9689 => x"384252e4",
     9690 => x"f80026a8",  9691 => x"5c200005",  9692 => x"fbffe884",
     9693 => x"78010001",  9694 => x"3821616c",  9695 => x"58200000",
     9696 => x"78010001",  9697 => x"3821616c",  9698 => x"28210000",
     9699 => x"78020001",  9700 => x"384252d8",  9701 => x"44200003",
     9702 => x"78020001",  9703 => x"384252d4",  9704 => x"78010001",
     9705 => x"382152ec",  9706 => x"f8000c05",  9707 => x"34010000",
     9708 => x"2b9d0004",  9709 => x"2b8b0008",  9710 => x"379c0008",
     9711 => x"c3a00000",  9712 => x"379cfff8",  9713 => x"5b8b0008",
     9714 => x"5b9d0004",  9715 => x"b8205800",  9716 => x"28210000",
     9717 => x"78020001",  9718 => x"384251f8",  9719 => x"f800268b",
     9720 => x"5c200003",  9721 => x"f80013c7",  9722 => x"e000000f",
     9723 => x"29610000",  9724 => x"78020001",  9725 => x"38425308",
     9726 => x"f8002684",  9727 => x"5c200003",  9728 => x"f80013c9",
     9729 => x"e0000008",  9730 => x"29610000",  9731 => x"78020001",
     9732 => x"3842530c",  9733 => x"f800267d",  9734 => x"3402ffea",
     9735 => x"5c200003",  9736 => x"f80013c7",  9737 => x"34020000",
     9738 => x"b8400800",  9739 => x"2b9d0004",  9740 => x"2b8b0008",
     9741 => x"379c0008",  9742 => x"c3a00000",  9743 => x"379cffec",
     9744 => x"5b8b0010",  9745 => x"5b8c000c",  9746 => x"5b8d0008",
     9747 => x"5b9d0004",  9748 => x"340b0000",  9749 => x"b8406800",
     9750 => x"340c0004",  9751 => x"37820014",  9752 => x"fbfffbd0",
     9753 => x"2b830014",  9754 => x"b5ab1000",  9755 => x"356b0001",
     9756 => x"30430000",  9757 => x"40220000",  9758 => x"6442002e",
     9759 => x"b4220800",  9760 => x"5d6cfff7",  9761 => x"2b9d0004",
     9762 => x"2b8b0010",  9763 => x"2b8c000c",  9764 => x"2b8d0008",
     9765 => x"379c0014",  9766 => x"c3a00000",  9767 => x"379cfff8",
     9768 => x"5b8b0008",  9769 => x"5b9d0004",  9770 => x"b8403000",
     9771 => x"40c30000",  9772 => x"40c40001",  9773 => x"40c50002",
     9774 => x"40c60003",  9775 => x"78020001",  9776 => x"38425318",
     9777 => x"b8205800",  9778 => x"f8000baf",  9779 => x"b9600800",
     9780 => x"2b9d0004",  9781 => x"2b8b0008",  9782 => x"379c0008",
     9783 => x"c3a00000",  9784 => x"379cffe0",  9785 => x"5b8b0008",
     9786 => x"5b9d0004",  9787 => x"b8205800",  9788 => x"28210000",
     9789 => x"44200005",  9790 => x"78020001",  9791 => x"38425004",
     9792 => x"f8002642",  9793 => x"5c200004",  9794 => x"37810020",
     9795 => x"f800050c",  9796 => x"e0000012",  9797 => x"29610000",
     9798 => x"78020001",  9799 => x"38425010",  9800 => x"f800263a",
     9801 => x"b8201800",  9802 => x"3402ffea",  9803 => x"5c200024",
     9804 => x"29610004",  9805 => x"44230022",  9806 => x"78020001",
     9807 => x"38427d90",  9808 => x"34030002",  9809 => x"58430000",
     9810 => x"37820020",  9811 => x"fbffffbc",  9812 => x"37810020",
     9813 => x"f8000503",  9814 => x"378b000c",  9815 => x"37820020",
     9816 => x"b9600800",  9817 => x"fbffffce",  9818 => x"78010001",
     9819 => x"38217d90",  9820 => x"28210000",  9821 => x"34020001",
     9822 => x"44220009",  9823 => x"44200004",  9824 => x"34020002",
     9825 => x"5c22000d",  9826 => x"e0000008",  9827 => x"78010001",
     9828 => x"38215324",  9829 => x"f8000b8a",  9830 => x"e0000008",
     9831 => x"78010001",  9832 => x"38215340",  9833 => x"e0000003",
     9834 => x"78010001",  9835 => x"38215360",  9836 => x"b9601000",
     9837 => x"f8000b82",  9838 => x"34020000",  9839 => x"b8400800",
     9840 => x"2b9d0004",  9841 => x"2b8b0008",  9842 => x"379c0020",
     9843 => x"c3a00000",  9844 => x"379cfffc",  9845 => x"5b9d0004",
     9846 => x"28210000",  9847 => x"44200005",  9848 => x"fbffdc00",
     9849 => x"78020001",  9850 => x"3842758c",  9851 => x"58410000",
     9852 => x"78020001",  9853 => x"3842758c",  9854 => x"28420000",
     9855 => x"78010001",  9856 => x"38215388",  9857 => x"f8000b6e",
     9858 => x"34010000",  9859 => x"2b9d0004",  9860 => x"379c0004",
     9861 => x"c3a00000",  9862 => x"379cfff0",  9863 => x"5b8b0008",
     9864 => x"5b9d0004",  9865 => x"b8205800",  9866 => x"28210000",
     9867 => x"5c200005",  9868 => x"78010001",  9869 => x"382153a8",
     9870 => x"f8000b61",  9871 => x"e0000010",  9872 => x"37820010",
     9873 => x"fbfffb3c",  9874 => x"29610004",  9875 => x"44200007",
     9876 => x"3782000c",  9877 => x"fbfffb38",  9878 => x"2b82000c",
     9879 => x"2b810010",  9880 => x"58220000",  9881 => x"e0000006",
     9882 => x"2b820010",  9883 => x"78010001",  9884 => x"382153d4",
     9885 => x"28430000",  9886 => x"f8000b51",  9887 => x"34010000",
     9888 => x"2b9d0004",  9889 => x"2b8b0008",  9890 => x"379c0010",
     9891 => x"c3a00000",  9892 => x"379cffe4",  9893 => x"5b8b0014",
     9894 => x"5b8c0010",  9895 => x"5b8d000c",  9896 => x"5b8e0008",
     9897 => x"5b9d0004",  9898 => x"b8205800",  9899 => x"78010001",
     9900 => x"38216178",  9901 => x"282e0014",  9902 => x"29610000",
     9903 => x"44200007",  9904 => x"29620004",  9905 => x"5c400005",
     9906 => x"78010001",  9907 => x"382153e4",  9908 => x"f8000b3b",
     9909 => x"e000001a",  9910 => x"29620004",  9911 => x"780d0001",
     9912 => x"780c0001",  9913 => x"39ad8ec8",  9914 => x"398c8ecc",
     9915 => x"4440000f",  9916 => x"3782001c",  9917 => x"fbfffb2b",
     9918 => x"29610004",  9919 => x"37820018",  9920 => x"fbfffb28",
     9921 => x"2b81001c",  9922 => x"2b8b0018",  9923 => x"59c10018",
     9924 => x"59a10000",  9925 => x"598b0000",  9926 => x"f8000c9a",
     9927 => x"b42b0800",  9928 => x"59c1001c",  9929 => x"e0000006",
     9930 => x"29a20000",  9931 => x"29830000",  9932 => x"78010001",
     9933 => x"38215414",  9934 => x"f8000b21",  9935 => x"34010000",
     9936 => x"2b9d0004",  9937 => x"2b8b0014",  9938 => x"2b8c0010",
     9939 => x"2b8d000c",  9940 => x"2b8e0008",  9941 => x"379c001c",
     9942 => x"c3a00000",  9943 => x"379cfff4",  9944 => x"5b8b000c",
     9945 => x"5b8c0008",  9946 => x"5b9d0004",  9947 => x"b8205800",
     9948 => x"28210000",  9949 => x"4420000b",  9950 => x"78020001",
     9951 => x"384250e0",  9952 => x"f80025a2",  9953 => x"b8206000",
     9954 => x"5c200006",  9955 => x"f8001670",  9956 => x"4c2c0025",
     9957 => x"78010001",  9958 => x"38215438",  9959 => x"e000000e",
     9960 => x"29610004",  9961 => x"44200011",  9962 => x"29610000",
     9963 => x"78020001",  9964 => x"384250fc",  9965 => x"f8002595",
     9966 => x"b8206000",  9967 => x"5c20000b",  9968 => x"b9600800",
     9969 => x"f8001677",  9970 => x"4c2c0005",  9971 => x"78010001",
     9972 => x"38215458",  9973 => x"f8000afa",  9974 => x"e0000013",
     9975 => x"78010001",  9976 => x"38215474",  9977 => x"e3fffffc",
     9978 => x"29610000",  9979 => x"44200007",  9980 => x"78020001",
     9981 => x"38425148",  9982 => x"f8002584",  9983 => x"5c200003",
     9984 => x"f80016e2",  9985 => x"e0000008",  9986 => x"29610000",
     9987 => x"44200006",  9988 => x"78020001",  9989 => x"3842547c",
     9990 => x"f800257c",  9991 => x"5c200002",  9992 => x"fbfffaed",
     9993 => x"34010000",  9994 => x"2b9d0004",  9995 => x"2b8b000c",
     9996 => x"2b8c0008",  9997 => x"379c000c",  9998 => x"c3a00000",
     9999 => x"379cffd0", 10000 => x"5b8b0030", 10001 => x"5b8c002c",
    10002 => x"5b8d0028", 10003 => x"5b8e0024", 10004 => x"5b8f0020",
    10005 => x"5b90001c", 10006 => x"5b910018", 10007 => x"5b920014",
    10008 => x"5b930010", 10009 => x"5b94000c", 10010 => x"5b9d0008",
    10011 => x"b8609000", 10012 => x"78030001", 10013 => x"38635a60",
    10014 => x"b8406000", 10015 => x"b8400800", 10016 => x"28620000",
    10017 => x"f8002451", 10018 => x"78030001", 10019 => x"38635a60",
    10020 => x"28620000", 10021 => x"b8205800", 10022 => x"b9800800",
    10023 => x"f800243b", 10024 => x"b820a000", 10025 => x"3402003c",
    10026 => x"b9600800", 10027 => x"f8002447", 10028 => x"34020e10",
    10029 => x"b8207800", 10030 => x"b9600800", 10031 => x"f8002443",
    10032 => x"3402003c", 10033 => x"f8002431", 10034 => x"b8208000",
    10035 => x"34020e10", 10036 => x"b9600800", 10037 => x"f800242d",
    10038 => x"b8208800", 10039 => x"ba807000", 10040 => x"340b07b2",
    10041 => x"e000000f", 10042 => x"3402016d", 10043 => x"5d80000b",
    10044 => x"34020064", 10045 => x"b9600800", 10046 => x"f8002404",
    10047 => x"3402016e", 10048 => x"5c2c0006", 10049 => x"34020190",
    10050 => x"b9600800", 10051 => x"f80023ff", 10052 => x"64220000",
    10053 => x"3442016d", 10054 => x"c9c27000", 10055 => x"356b0001",
    10056 => x"216c0003", 10057 => x"3402016d", 10058 => x"5d80000b",
    10059 => x"34020064", 10060 => x"b9600800", 10061 => x"f80023f5",
    10062 => x"3402016e", 10063 => x"5c2c0006", 10064 => x"34020190",
    10065 => x"b9600800", 10066 => x"f80023f0", 10067 => x"64220000",
    10068 => x"3442016d", 10069 => x"51c2ffe5", 10070 => x"34020064",
    10071 => x"b9600800", 10072 => x"f80023ea", 10073 => x"34020190",
    10074 => x"b8209800", 10075 => x"b9600800", 10076 => x"f80023e6",
    10077 => x"78020001", 10078 => x"340d0000", 10079 => x"64250000",
    10080 => x"38425d48", 10081 => x"e000000d", 10082 => x"34040000",
    10083 => x"5d800004", 10084 => x"34040001", 10085 => x"5e6c0002",
    10086 => x"b8a02000", 10087 => x"0884000c", 10088 => x"b48d2000",
    10089 => x"3c840002", 10090 => x"35ad0001", 10091 => x"b4442000",
    10092 => x"28810000", 10093 => x"c9c17000", 10094 => x"34040000",
    10095 => x"5d800004", 10096 => x"34040001", 10097 => x"5e6c0002",
    10098 => x"b8a02000", 10099 => x"0884000c", 10100 => x"b48d2000",
    10101 => x"3c840002", 10102 => x"b4442000", 10103 => x"28810000",
    10104 => x"51c1ffea", 10105 => x"34010001", 10106 => x"35ce0001",
    10107 => x"4641001d", 10108 => x"780c0001", 10109 => x"34010002",
    10110 => x"398c7b2c", 10111 => x"46410028", 10112 => x"36810004",
    10113 => x"34020007", 10114 => x"f80023f0", 10115 => x"3c210002",
    10116 => x"78130001", 10117 => x"78020001", 10118 => x"3dad0002",
    10119 => x"38425dc4", 10120 => x"3a735da8", 10121 => x"b6619800",
    10122 => x"b44d6800", 10123 => x"78120001", 10124 => x"2a630000",
    10125 => x"29a40000", 10126 => x"3a525484", 10127 => x"b9800800",
    10128 => x"ba401000", 10129 => x"b9c02800", 10130 => x"b9603000",
    10131 => x"ba203800", 10132 => x"ba004000", 10133 => x"5b8f0004",
    10134 => x"f8000a4b", 10135 => x"e000001a", 10136 => x"78010001",
    10137 => x"3dad0002", 10138 => x"38215dc4", 10139 => x"b42d6800",
    10140 => x"29a30000", 10141 => x"78010001", 10142 => x"78020001",
    10143 => x"384254a4", 10144 => x"b9c02000", 10145 => x"ba202800",
    10146 => x"ba003000", 10147 => x"b9e03800", 10148 => x"38217b2c",
    10149 => x"f8000a3c", 10150 => x"e000000b", 10151 => x"78020001",
    10152 => x"b9800800", 10153 => x"384254bc", 10154 => x"b9601800",
    10155 => x"35a40001", 10156 => x"b9c02800", 10157 => x"ba203000",
    10158 => x"ba003800", 10159 => x"b9e04000", 10160 => x"f8000a31",
    10161 => x"78010001", 10162 => x"38217b2c", 10163 => x"2b9d0008",
    10164 => x"2b8b0030", 10165 => x"2b8c002c", 10166 => x"2b8d0028",
    10167 => x"2b8e0024", 10168 => x"2b8f0020", 10169 => x"2b90001c",
    10170 => x"2b910018", 10171 => x"2b920014", 10172 => x"2b930010",
    10173 => x"2b94000c", 10174 => x"379c0030", 10175 => x"c3a00000",
    10176 => x"379cffdc", 10177 => x"5b8b0008", 10178 => x"5b9d0004",
    10179 => x"5b840014", 10180 => x"20240080", 10181 => x"64840000",
    10182 => x"5b830010", 10183 => x"78030001", 10184 => x"b8204800",
    10185 => x"b8600800", 10186 => x"34030002", 10187 => x"5b82000c",
    10188 => x"b8405800", 10189 => x"382154dc", 10190 => x"c8641000",
    10191 => x"2123007f", 10192 => x"5b850018", 10193 => x"5b86001c",
    10194 => x"5b870020", 10195 => x"5b880024", 10196 => x"f8000a1b",
    10197 => x"37820010", 10198 => x"b9600800", 10199 => x"f80009f6",
    10200 => x"78010001", 10201 => x"382154e8", 10202 => x"f8000a15",
    10203 => x"2b9d0004", 10204 => x"2b8b0008", 10205 => x"379c0024",
    10206 => x"c3a00000", 10207 => x"379cffe0", 10208 => x"5b8b000c",
    10209 => x"5b8c0008", 10210 => x"5b9d0004", 10211 => x"b8404800",
    10212 => x"78020001", 10213 => x"b8205000", 10214 => x"b8400800",
    10215 => x"b8605800", 10216 => x"b9401000", 10217 => x"b9201800",
    10218 => x"382154ec", 10219 => x"b8806000", 10220 => x"5b840010",
    10221 => x"5b850014", 10222 => x"5b860018", 10223 => x"5b87001c",
    10224 => x"5b880020", 10225 => x"f80009fe", 10226 => x"21620080",
    10227 => x"78030001", 10228 => x"64420000", 10229 => x"b8600800",
    10230 => x"34030002", 10231 => x"c8621000", 10232 => x"382154dc",
    10233 => x"2163007f", 10234 => x"f80009f5", 10235 => x"37820014",
    10236 => x"b9800800", 10237 => x"f80009d0", 10238 => x"78010001",
    10239 => x"382154e8", 10240 => x"f80009ef", 10241 => x"2b9d0004",
    10242 => x"2b8b000c", 10243 => x"2b8c0008", 10244 => x"379c0020",
    10245 => x"c3a00000", 10246 => x"379cfffc", 10247 => x"5b9d0004",
    10248 => x"78010001", 10249 => x"382154f8", 10250 => x"f80009e5",
    10251 => x"2b9d0004", 10252 => x"379c0004", 10253 => x"c3a00000",
    10254 => x"40240000", 10255 => x"3402002d", 10256 => x"34030001",
    10257 => x"5c820003", 10258 => x"34210001", 10259 => x"3403ffff",
    10260 => x"34020000", 10261 => x"34050009", 10262 => x"e0000004",
    10263 => x"0842000a", 10264 => x"34210001", 10265 => x"b4821000",
    10266 => x"40240000", 10267 => x"3484ffd0", 10268 => x"208600ff",
    10269 => x"50a6fffa", 10270 => x"88430800", 10271 => x"c3a00000",
    10272 => x"379cfff4", 10273 => x"5b8b000c", 10274 => x"5b8c0008",
    10275 => x"5b9d0004", 10276 => x"b8206000", 10277 => x"f8000f8a",
    10278 => x"342b0001", 10279 => x"f8000f88", 10280 => x"5c2bffff",
    10281 => x"b9800800", 10282 => x"e0000002", 10283 => x"3421ffff",
    10284 => x"4820ffff", 10285 => x"f8000f82", 10286 => x"c82b0800",
    10287 => x"2b9d0004", 10288 => x"2b8b000c", 10289 => x"2b8c0008",
    10290 => x"379c000c", 10291 => x"c3a00000", 10292 => x"379cfff0",
    10293 => x"5b8b0010", 10294 => x"5b8c000c", 10295 => x"5b8d0008",
    10296 => x"5b9d0004", 10297 => x"340b0400", 10298 => x"340c0400",
    10299 => x"e0000003", 10300 => x"b58b6000", 10301 => x"3d6b0001",
    10302 => x"b9800800", 10303 => x"fbffffe1", 10304 => x"4420fffc",
    10305 => x"158c0001", 10306 => x"156b0002", 10307 => x"e0000009",
    10308 => x"b56c6800", 10309 => x"b9a00800", 10310 => x"fbffffda",
    10311 => x"5c200002", 10312 => x"b9a06000", 10313 => x"0161001f",
    10314 => x"b42b5800", 10315 => x"156b0001", 10316 => x"5d60fff8",
    10317 => x"78010001", 10318 => x"38217b6c", 10319 => x"582c0000",
    10320 => x"78010001", 10321 => x"b9801000", 10322 => x"38215550",
    10323 => x"f800099c", 10324 => x"2b9d0004", 10325 => x"2b8b0010",
    10326 => x"2b8c000c", 10327 => x"2b8d0008", 10328 => x"379c0010",
    10329 => x"c3a00000", 10330 => x"379cfffc", 10331 => x"5b9d0004",
    10332 => x"78020001", 10333 => x"38427b6c", 10334 => x"28430000",
    10335 => x"34042710", 10336 => x"0865000a", 10337 => x"e0000004",
    10338 => x"3442ffff", 10339 => x"4840ffff", 10340 => x"3421d8f0",
    10341 => x"50810003", 10342 => x"b8a01000", 10343 => x"e3fffffc",
    10344 => x"88230800", 10345 => x"340203e8", 10346 => x"f80022f8",
    10347 => x"e0000002", 10348 => x"3421ffff", 10349 => x"4820ffff",
    10350 => x"34010000", 10351 => x"2b9d0004", 10352 => x"379c0004",
    10353 => x"c3a00000", 10354 => x"b8202800", 10355 => x"5c800002",
    10356 => x"b8602000", 10357 => x"b8803000", 10358 => x"50640002",
    10359 => x"b8603000", 10360 => x"b4260800", 10361 => x"e000000e",
    10362 => x"2c460002", 10363 => x"2847000c", 10364 => x"b4e63800",
    10365 => x"40e60000", 10366 => x"30a60000", 10367 => x"2c470002",
    10368 => x"2c460006", 10369 => x"34a50001", 10370 => x"34e70001",
    10371 => x"20e7ffff", 10372 => x"0c470002", 10373 => x"5cc70002",
    10374 => x"0c400002", 10375 => x"5ca1fff3", 10376 => x"5083000b",
    10377 => x"2c410002", 10378 => x"b4610800", 10379 => x"c8242000",
    10380 => x"0c440002", 10381 => x"2c410006", 10382 => x"e0000003",
    10383 => x"c8812000", 10384 => x"0c440002", 10385 => x"2c440002",
    10386 => x"5481fffd", 10387 => x"b8600800", 10388 => x"c3a00000",
    10389 => x"b4432800", 10390 => x"e000000d", 10391 => x"2c240000",
    10392 => x"2826000c", 10393 => x"40470000", 10394 => x"34420001",
    10395 => x"b4c43000", 10396 => x"30c70000", 10397 => x"34840001",
    10398 => x"2c260006", 10399 => x"2084ffff", 10400 => x"0c240000",
    10401 => x"5cc40002", 10402 => x"0c200000", 10403 => x"5c45fff4",
    10404 => x"b8600800", 10405 => x"c3a00000", 10406 => x"379cffc8",
    10407 => x"5b8b001c", 10408 => x"5b8c0018", 10409 => x"5b8d0014",
    10410 => x"5b8e0010", 10411 => x"5b8f000c", 10412 => x"5b900008",
    10413 => x"5b9d0004", 10414 => x"780b0001", 10415 => x"780c0001",
    10416 => x"396b7d80", 10417 => x"398c7ba0", 10418 => x"b9600800",
    10419 => x"b9801000", 10420 => x"340301e0", 10421 => x"37840020",
    10422 => x"f8000d94", 10423 => x"b8206800", 10424 => x"340f0000",
    10425 => x"4c010061", 10426 => x"2d62000c", 10427 => x"0f800038",
    10428 => x"38018100", 10429 => x"5c41000e", 10430 => x"b9801000",
    10431 => x"34030002", 10432 => x"37810038", 10433 => x"f8002302",
    10434 => x"78010001", 10435 => x"78020001", 10436 => x"38217d8c",
    10437 => x"38427ba2", 10438 => x"34030002", 10439 => x"780c0001",
    10440 => x"f80022fb", 10441 => x"35adfffc", 10442 => x"398c7ba4",
    10443 => x"78010001", 10444 => x"2f820038", 10445 => x"3821757c",
    10446 => x"28210000", 10447 => x"20420fff", 10448 => x"340f0000",
    10449 => x"5c410049", 10450 => x"41820000", 10451 => x"34010045",
    10452 => x"34030000", 10453 => x"5c410008", 10454 => x"41820009",
    10455 => x"34010011", 10456 => x"5c410005", 10457 => x"41830016",
    10458 => x"41810017", 10459 => x"3c630008", 10460 => x"b8611800",
    10461 => x"78010001", 10462 => x"78020001", 10463 => x"38217d80",
    10464 => x"38427b70", 10465 => x"2c27000c", 10466 => x"34460030",
    10467 => x"34040000", 10468 => x"340b0000", 10469 => x"e000000c",
    10470 => x"28410000", 10471 => x"44200009", 10472 => x"2c25000c",
    10473 => x"5ca70007", 10474 => x"2c25000e", 10475 => x"5c600003",
    10476 => x"44a30038", 10477 => x"e0000003", 10478 => x"5ca30002",
    10479 => x"b8202000", 10480 => x"34420004", 10481 => x"5c46fff5",
    10482 => x"44800002", 10483 => x"b8805800", 10484 => x"340f0001",
    10485 => x"45600025", 10486 => x"2d700028", 10487 => x"35a10028",
    10488 => x"48300022", 10489 => x"356e0024", 10490 => x"3782003a",
    10491 => x"34030002", 10492 => x"b9c00800", 10493 => x"0f8d003a",
    10494 => x"fbffff97", 10495 => x"ca016800", 10496 => x"21adffff",
    10497 => x"0d6d0028", 10498 => x"37820020", 10499 => x"34030018",
    10500 => x"b9c00800", 10501 => x"fbffff90", 10502 => x"c9a16800",
    10503 => x"21adffff", 10504 => x"78020001", 10505 => x"0d6d0028",
    10506 => x"38427d80", 10507 => x"3403000e", 10508 => x"b9c00800",
    10509 => x"fbffff88", 10510 => x"c9a16800", 10511 => x"2f83003a",
    10512 => x"21adffff", 10513 => x"0d6d0028", 10514 => x"b9c00800",
    10515 => x"b9801000", 10516 => x"fbffff81", 10517 => x"c9a10800",
    10518 => x"0d610028", 10519 => x"2d61002c", 10520 => x"34210001",
    10521 => x"0d61002c", 10522 => x"b9e00800", 10523 => x"2b9d0004",
    10524 => x"2b8b001c", 10525 => x"2b8c0018", 10526 => x"2b8d0014",
    10527 => x"2b8e0010", 10528 => x"2b8f000c", 10529 => x"2b900008",
    10530 => x"379c0038", 10531 => x"c3a00000", 10532 => x"b8205800",
    10533 => x"e3ffffcb", 10534 => x"379cfffc", 10535 => x"5b9d0004",
    10536 => x"b8400800", 10537 => x"f80009ce", 10538 => x"34010000",
    10539 => x"2b9d0004", 10540 => x"379c0004", 10541 => x"c3a00000",
    10542 => x"78020001", 10543 => x"38427b70", 10544 => x"34430030",
    10545 => x"e0000004", 10546 => x"28440000", 10547 => x"34420004",
    10548 => x"5881001c", 10549 => x"5c43fffd", 10550 => x"c3a00000",
    10551 => x"379cff24", 10552 => x"5b8b0014", 10553 => x"5b8c0010",
    10554 => x"5b8d000c", 10555 => x"5b8e0008", 10556 => x"5b9d0004",
    10557 => x"78050001", 10558 => x"b8205800", 10559 => x"b8406000",
    10560 => x"b8607000", 10561 => x"b8806800", 10562 => x"38a57b70",
    10563 => x"34010000", 10564 => x"3402000c", 10565 => x"28a30000",
    10566 => x"34a50004", 10567 => x"5c600009", 10568 => x"3c220002",
    10569 => x"78050001", 10570 => x"38a57b70", 10571 => x"b4a22800",
    10572 => x"58ab0000", 10573 => x"3402000c", 10574 => x"5c22000a",
    10575 => x"e0000003", 10576 => x"34210001", 10577 => x"5c22fff4",
    10578 => x"78010001", 10579 => x"78020001", 10580 => x"38425df4",
    10581 => x"38215568", 10582 => x"f8000899", 10583 => x"e0000020",
    10584 => x"78020001", 10585 => x"37810018", 10586 => x"38425584",
    10587 => x"fbfff70a", 10588 => x"4801001b", 10589 => x"b9600800",
    10590 => x"34020000", 10591 => x"34030012", 10592 => x"f80022e1",
    10593 => x"45800005", 10594 => x"b9600800", 10595 => x"b9801000",
    10596 => x"34030012", 10597 => x"f800225e", 10598 => x"0d60000e",
    10599 => x"5dc00004", 10600 => x"34010800", 10601 => x"0d61000c",
    10602 => x"0d6d000e", 10603 => x"35610012", 10604 => x"f800098b",
    10605 => x"2b8100d0", 10606 => x"0d600026", 10607 => x"0d600024",
    10608 => x"5961001c", 10609 => x"2b8100b8", 10610 => x"0d60002c",
    10611 => x"59610020", 10612 => x"2d61002a", 10613 => x"0d610028",
    10614 => x"e0000002", 10615 => x"340b0000", 10616 => x"b9600800",
    10617 => x"2b9d0004", 10618 => x"2b8b0014", 10619 => x"2b8c0010",
    10620 => x"2b8d000c", 10621 => x"2b8e0008", 10622 => x"379c00dc",
    10623 => x"c3a00000", 10624 => x"78020001", 10625 => x"38427b70",
    10626 => x"34430030", 10627 => x"e0000005", 10628 => x"28440000",
    10629 => x"5c810002", 10630 => x"58400000", 10631 => x"34420004",
    10632 => x"5c43fffc", 10633 => x"34010000", 10634 => x"c3a00000",
    10635 => x"379cffe8", 10636 => x"5b8b0018", 10637 => x"5b8c0014",
    10638 => x"5b8d0010", 10639 => x"5b8e000c", 10640 => x"5b8f0008",
    10641 => x"5b9d0004", 10642 => x"b8205800", 10643 => x"59620010",
    10644 => x"b8407000", 10645 => x"b8807800", 10646 => x"b8a06000",
    10647 => x"282d0008", 10648 => x"44600005", 10649 => x"b8a00800",
    10650 => x"3402fc18", 10651 => x"f800217a", 10652 => x"b42d6800",
    10653 => x"c9cf2000", 10654 => x"b8801800", 10655 => x"4c800002",
    10656 => x"b48c1800", 10657 => x"0181001f", 10658 => x"b42c0800",
    10659 => x"14210001", 10660 => x"b4242000", 10661 => x"4c800002",
    10662 => x"b48c2000", 10663 => x"49840002", 10664 => x"c88c2000",
    10665 => x"09820003", 10666 => x"1445001f", 10667 => x"00a5001e",
    10668 => x"b4a21000", 10669 => x"14420002", 10670 => x"48620006",
    10671 => x"1582001f", 10672 => x"0042001e", 10673 => x"b44c1000",
    10674 => x"14420002", 10675 => x"4c62000d", 10676 => x"b4812000",
    10677 => x"596d0008", 10678 => x"5964000c", 10679 => x"4984000a",
    10680 => x"c88c2000", 10681 => x"5964000c", 10682 => x"b9800800",
    10683 => x"340203e8", 10684 => x"f8002159", 10685 => x"b5a10800",
    10686 => x"59610008", 10687 => x"e0000002", 10688 => x"5963000c",
    10689 => x"78030001", 10690 => x"38635a3c", 10691 => x"29610008",
    10692 => x"28620000", 10693 => x"4c41000d", 10694 => x"78030001",
    10695 => x"38635a40", 10696 => x"28620000", 10697 => x"29630000",
    10698 => x"b4220800", 10699 => x"29620004", 10700 => x"59610008",
    10701 => x"34410001", 10702 => x"f4411000", 10703 => x"59610004",
    10704 => x"b4431000", 10705 => x"59620000", 10706 => x"2b9d0004",
    10707 => x"2b8b0018", 10708 => x"2b8c0014", 10709 => x"2b8d0010",
    10710 => x"2b8e000c", 10711 => x"2b8f0008", 10712 => x"379c0018",
    10713 => x"c3a00000", 10714 => x"379cffb4", 10715 => x"5b8b0024",
    10716 => x"5b8c0020", 10717 => x"5b8d001c", 10718 => x"5b8e0018",
    10719 => x"5b8f0014", 10720 => x"5b900010", 10721 => x"5b91000c",
    10722 => x"5b920008", 10723 => x"5b9d0004", 10724 => x"b8406800",
    10725 => x"2c22002c", 10726 => x"b8a05800", 10727 => x"b8206000",
    10728 => x"b8609000", 10729 => x"b8807800", 10730 => x"34050000",
    10731 => x"44400055", 10732 => x"342e0024", 10733 => x"2c310028",
    10734 => x"3442ffff", 10735 => x"0c22002c", 10736 => x"34030002",
    10737 => x"b9c01000", 10738 => x"34040000", 10739 => x"3781004e",
    10740 => x"fbfffe7e", 10741 => x"b6218800", 10742 => x"2231ffff",
    10743 => x"0d910028", 10744 => x"b9c01000", 10745 => x"34030018",
    10746 => x"34040000", 10747 => x"37810028", 10748 => x"fbfffe76",
    10749 => x"b6218800", 10750 => x"2231ffff", 10751 => x"37900040",
    10752 => x"0d910028", 10753 => x"b9c01000", 10754 => x"3403000e",
    10755 => x"34040000", 10756 => x"ba000800", 10757 => x"fbfffe6d",
    10758 => x"b6218800", 10759 => x"2f83004e", 10760 => x"2231ffff",
    10761 => x"b9c01000", 10762 => x"b9e02000", 10763 => x"0d910028",
    10764 => x"ba400800", 10765 => x"fbfffe65", 10766 => x"b6210800",
    10767 => x"0d810028", 10768 => x"2f81004c", 10769 => x"78030001",
    10770 => x"3863757c", 10771 => x"0da1000c", 10772 => x"28610000",
    10773 => x"37820046", 10774 => x"34030006", 10775 => x"0da10010",
    10776 => x"b9a00800", 10777 => x"f80021aa", 10778 => x"35a10006",
    10779 => x"ba001000", 10780 => x"34030006", 10781 => x"f80021a6",
    10782 => x"4560001e", 10783 => x"2b810038", 10784 => x"59610014",
    10785 => x"2b81002c", 10786 => x"59610018", 10787 => x"34010000",
    10788 => x"f8001e87", 10789 => x"b8206800", 10790 => x"35620010",
    10791 => x"34030000", 10792 => x"34010000", 10793 => x"f8001e2d",
    10794 => x"2b810030", 10795 => x"43820028", 10796 => x"2b83002c",
    10797 => x"59610000", 10798 => x"2b810034", 10799 => x"2984001c",
    10800 => x"5960000c", 10801 => x"59610004", 10802 => x"2b810038",
    10803 => x"34051f40", 10804 => x"59610008", 10805 => x"21a100ff",
    10806 => x"64210000", 10807 => x"a0220800", 10808 => x"29620010",
    10809 => x"5961001c", 10810 => x"b9600800", 10811 => x"fbffff50",
    10812 => x"2f81004e", 10813 => x"b9e02800", 10814 => x"502f0002",
    10815 => x"b8202800", 10816 => x"b8a00800", 10817 => x"2b9d0004",
    10818 => x"2b8b0024", 10819 => x"2b8c0020", 10820 => x"2b8d001c",
    10821 => x"2b8e0018", 10822 => x"2b8f0014", 10823 => x"2b900010",
    10824 => x"2b91000c", 10825 => x"2b920008", 10826 => x"379c004c",
    10827 => x"c3a00000", 10828 => x"379cffc0", 10829 => x"5b8b0014",
    10830 => x"5b8c0010", 10831 => x"5b8d000c", 10832 => x"5b8e0008",
    10833 => x"5b9d0004", 10834 => x"b8206000", 10835 => x"b8607000",
    10836 => x"37810030", 10837 => x"34030006", 10838 => x"b8a05800",
    10839 => x"b8806800", 10840 => x"f800216b", 10841 => x"37810036",
    10842 => x"35820012", 10843 => x"34030006", 10844 => x"f8002167",
    10845 => x"78010001", 10846 => x"3821757c", 10847 => x"28250000",
    10848 => x"2d81000c", 10849 => x"44a00009", 10850 => x"34028100",
    10851 => x"0f82003c", 10852 => x"2d820018", 10853 => x"0f810040",
    10854 => x"3c42000d", 10855 => x"b8452800", 10856 => x"0f85003e",
    10857 => x"e0000002", 10858 => x"0f81003c", 10859 => x"37810030",
    10860 => x"b9c01000", 10861 => x"b9a01800", 10862 => x"37840018",
    10863 => x"f8000c86", 10864 => x"4560000a", 10865 => x"2b820020",
    10866 => x"5960000c", 10867 => x"59620000", 10868 => x"2b820024",
    10869 => x"59620004", 10870 => x"2b820028", 10871 => x"59620008",
    10872 => x"43820018", 10873 => x"5962001c", 10874 => x"2b9d0004",
    10875 => x"2b8b0014", 10876 => x"2b8c0010", 10877 => x"2b8d000c",
    10878 => x"2b8e0008", 10879 => x"379c0040", 10880 => x"c3a00000",
    10881 => x"c3a00000", 10882 => x"379cffe4", 10883 => x"5b8b0008",
    10884 => x"5b9d0004", 10885 => x"78010001", 10886 => x"34020000",
    10887 => x"34030000", 10888 => x"34040044", 10889 => x"38216874",
    10890 => x"fbfffead", 10891 => x"78020001", 10892 => x"38427d94",
    10893 => x"58410000", 10894 => x"78010001", 10895 => x"34040025",
    10896 => x"34020000", 10897 => x"34030000", 10898 => x"382168a8",
    10899 => x"fbfffea4", 10900 => x"78020001", 10901 => x"378b000c",
    10902 => x"38427da4", 10903 => x"58410000", 10904 => x"34030012",
    10905 => x"b9600800", 10906 => x"34020000", 10907 => x"f80021a6",
    10908 => x"34010800", 10909 => x"0f810018", 10910 => x"78010001",
    10911 => x"b9601000", 10912 => x"34030001", 10913 => x"34040000",
    10914 => x"382168dc", 10915 => x"fbfffe94", 10916 => x"78020001",
    10917 => x"38427da0", 10918 => x"58410000", 10919 => x"fbffffda",
    10920 => x"2b9d0004", 10921 => x"2b8b0008", 10922 => x"379c001c",
    10923 => x"c3a00000", 10924 => x"34010000", 10925 => x"c3a00000",
    10926 => x"379cfe34", 10927 => x"5b8b001c", 10928 => x"5b8c0018",
    10929 => x"5b8d0014", 10930 => x"5b8e0010", 10931 => x"5b8f000c",
    10932 => x"5b900008", 10933 => x"5b9d0004", 10934 => x"78010001",
    10935 => x"382192a0", 10936 => x"28220000", 10937 => x"34010001",
    10938 => x"5c410006", 10939 => x"78010001", 10940 => x"38217d90",
    10941 => x"28230000", 10942 => x"5c620002", 10943 => x"58200000",
    10944 => x"78020001", 10945 => x"38427d94", 10946 => x"28410000",
    10947 => x"378b0020", 10948 => x"378201b0", 10949 => x"34040190",
    10950 => x"b9601800", 10951 => x"34050000", 10952 => x"fbffff12",
    10953 => x"78040001", 10954 => x"38847d90", 10955 => x"b8201000",
    10956 => x"28810000", 10957 => x"340c0000", 10958 => x"5c200023",
    10959 => x"4c220003", 10960 => x"b9600800", 10961 => x"f800027a",
    10962 => x"f8000cdd", 10963 => x"78020001", 10964 => x"38427d98",
    10965 => x"28430000", 10966 => x"5c600003", 10967 => x"58410000",
    10968 => x"e0000006", 10969 => x"346303e8", 10970 => x"c8230800",
    10971 => x"340c0000", 10972 => x"48010015", 10973 => x"58430000",
    10974 => x"78010001", 10975 => x"38217d9c", 10976 => x"28230000",
    10977 => x"378c01b0", 10978 => x"378b0020", 10979 => x"34630001",
    10980 => x"58230000", 10981 => x"b9601000", 10982 => x"b9800800",
    10983 => x"f8000200", 10984 => x"78050001", 10985 => x"38a57d94",
    10986 => x"b8202000", 10987 => x"28a10000", 10988 => x"b9801000",
    10989 => x"b9601800", 10990 => x"34050000", 10991 => x"fbffff5d",
    10992 => x"340c0001", 10993 => x"780b0001", 10994 => x"396b7da0",
    10995 => x"29610000", 10996 => x"378e01b0", 10997 => x"378d0020",
    10998 => x"34040080", 10999 => x"b9c01000", 11000 => x"b9a01800",
    11001 => x"34050000", 11002 => x"fbfffee0", 11003 => x"b8202000",
    11004 => x"340f0000", 11005 => x"4c010010", 11006 => x"78030001",
    11007 => x"38637d90", 11008 => x"28610000", 11009 => x"4420000c",
    11010 => x"b8801000", 11011 => x"b9a00800", 11012 => x"f8000108",
    11013 => x"b8202000", 11014 => x"340f0001", 11015 => x"4c010006",
    11016 => x"29610000", 11017 => x"b9c01000", 11018 => x"b9a01800",
    11019 => x"34050000", 11020 => x"fbffff40", 11021 => x"780b0001",
    11022 => x"396b7da4", 11023 => x"29610000", 11024 => x"379001b0",
    11025 => x"378d0020", 11026 => x"ba001000", 11027 => x"b9a01800",
    11028 => x"34040020", 11029 => x"34050000", 11030 => x"fbfffec4",
    11031 => x"340e0000", 11032 => x"4c010019", 11033 => x"378101c4",
    11034 => x"34020000", 11035 => x"f8001030", 11036 => x"78020001",
    11037 => x"38425a64", 11038 => x"28410000", 11039 => x"2b8201c8",
    11040 => x"34030004", 11041 => x"340e0001", 11042 => x"b4410800",
    11043 => x"5b8101cc", 11044 => x"378201cc", 11045 => x"3781003c",
    11046 => x"f800209d", 11047 => x"b9a00800", 11048 => x"34020020",
    11049 => x"34030000", 11050 => x"f8000143", 11051 => x"29610000",
    11052 => x"ba001000", 11053 => x"b9a01800", 11054 => x"34040020",
    11055 => x"34050000", 11056 => x"fbffff1c", 11057 => x"fbffff7b",
    11058 => x"b5ec6000", 11059 => x"b5810800", 11060 => x"b42e7000",
    11061 => x"7dc10000", 11062 => x"2b9d0004", 11063 => x"2b8b001c",
    11064 => x"2b8c0018", 11065 => x"2b8d0014", 11066 => x"2b8e0010",
    11067 => x"2b8f000c", 11068 => x"2b900008", 11069 => x"379c01cc",
    11070 => x"c3a00000", 11071 => x"34030000", 11072 => x"34040000",
    11073 => x"e0000005", 11074 => x"2c250000", 11075 => x"34840001",
    11076 => x"34210002", 11077 => x"b4651800", 11078 => x"4844fffc",
    11079 => x"00610010", 11080 => x"2063ffff", 11081 => x"b4611800",
    11082 => x"00610010", 11083 => x"b4231800", 11084 => x"a4600800",
    11085 => x"2021ffff", 11086 => x"c3a00000", 11087 => x"379cfffc",
    11088 => x"5b9d0004", 11089 => x"78020001", 11090 => x"38427da8",
    11091 => x"34030004", 11092 => x"f800206f", 11093 => x"2b9d0004",
    11094 => x"379c0004", 11095 => x"c3a00000", 11096 => x"379cfff0",
    11097 => x"5b8b0010", 11098 => x"5b8c000c", 11099 => x"5b8d0008",
    11100 => x"5b9d0004", 11101 => x"78030001", 11102 => x"780b0001",
    11103 => x"396b7da8", 11104 => x"b8206000", 11105 => x"386392b8",
    11106 => x"286d0000", 11107 => x"b9600800", 11108 => x"b9801000",
    11109 => x"34030004", 11110 => x"f800205d", 11111 => x"41620000",
    11112 => x"41610001", 11113 => x"3c420018", 11114 => x"3c210010",
    11115 => x"b8411000", 11116 => x"41610003", 11117 => x"b8411000",
    11118 => x"41610002", 11119 => x"3c210008", 11120 => x"b8415800",
    11121 => x"29a10018", 11122 => x"b9800800", 11123 => x"f8000e81",
    11124 => x"5d600004", 11125 => x"78010001", 11126 => x"38217d90",
    11127 => x"58200000", 11128 => x"78010001", 11129 => x"38217d9c",
    11130 => x"58200000", 11131 => x"2b9d0004", 11132 => x"2b8b0010",
    11133 => x"2b8c000c", 11134 => x"2b8d0008", 11135 => x"379c0010",
    11136 => x"c3a00000", 11137 => x"379cfffc", 11138 => x"5b9d0004",
    11139 => x"b8201000", 11140 => x"3401ffff", 11141 => x"44400006",
    11142 => x"34410010", 11143 => x"78020001", 11144 => x"38427da8",
    11145 => x"34030004", 11146 => x"f8002018", 11147 => x"2b9d0004",
    11148 => x"379c0004", 11149 => x"c3a00000", 11150 => x"379cff34",
    11151 => x"5b8b0028", 11152 => x"5b8c0024", 11153 => x"5b8d0020",
    11154 => x"5b8e001c", 11155 => x"5b8f0018", 11156 => x"5b900014",
    11157 => x"5b910010", 11158 => x"5b92000c", 11159 => x"5b930008",
    11160 => x"5b9d0004", 11161 => x"78010001", 11162 => x"38217d90",
    11163 => x"28210000", 11164 => x"340b0000", 11165 => x"44200047",
    11166 => x"780c0001", 11167 => x"398c808c", 11168 => x"29810000",
    11169 => x"378f00ac", 11170 => x"378e002c", 11171 => x"b9e01000",
    11172 => x"b9c01800", 11173 => x"34040080", 11174 => x"34050000",
    11175 => x"fbfffe33", 11176 => x"4c01003c", 11177 => x"3402001b",
    11178 => x"340b0001", 11179 => x"4c410039", 11180 => x"378d00c8",
    11181 => x"b9a00800", 11182 => x"fbffffa1", 11183 => x"43810032",
    11184 => x"5c200034", 11185 => x"43810033", 11186 => x"5c2b0032",
    11187 => x"37900044", 11188 => x"ba000800", 11189 => x"b9a01000",
    11190 => x"34030004", 11191 => x"f8001feb", 11192 => x"5c20002c",
    11193 => x"379100c0", 11194 => x"37930034", 11195 => x"ba601000",
    11196 => x"34030006", 11197 => x"ba200800", 11198 => x"f8002005",
    11199 => x"3792003a", 11200 => x"ba401000", 11201 => x"34030004",
    11202 => x"378100cc", 11203 => x"f8002000", 11204 => x"34010008",
    11205 => x"3381002e", 11206 => x"34010006", 11207 => x"33810030",
    11208 => x"34010004", 11209 => x"33810031", 11210 => x"34010002",
    11211 => x"33810033", 11212 => x"ba600800", 11213 => x"3380002c",
    11214 => x"338b002d", 11215 => x"3380002f", 11216 => x"33800032",
    11217 => x"f8000726", 11218 => x"b9a01000", 11219 => x"34030004",
    11220 => x"ba400800", 11221 => x"f8001fee", 11222 => x"ba201000",
    11223 => x"34030006", 11224 => x"3781003e", 11225 => x"f8001fea",
    11226 => x"378200cc", 11227 => x"34030004", 11228 => x"ba000800",
    11229 => x"f8001fe6", 11230 => x"29810000", 11231 => x"b9e01000",
    11232 => x"b9c01800", 11233 => x"3404001c", 11234 => x"34050000",
    11235 => x"fbfffe69", 11236 => x"b9600800", 11237 => x"2b9d0004",
    11238 => x"2b8b0028", 11239 => x"2b8c0024", 11240 => x"2b8d0020",
    11241 => x"2b8e001c", 11242 => x"2b8f0018", 11243 => x"2b900014",
    11244 => x"2b910010", 11245 => x"2b92000c", 11246 => x"2b930008",
    11247 => x"379c00cc", 11248 => x"c3a00000", 11249 => x"379cffe4",
    11250 => x"5b8b0008", 11251 => x"5b9d0004", 11252 => x"378b000c",
    11253 => x"b9600800", 11254 => x"34020000", 11255 => x"34030012",
    11256 => x"f8002049", 11257 => x"b9600800", 11258 => x"340200ff",
    11259 => x"34030006", 11260 => x"f8002045", 11261 => x"34010806",
    11262 => x"0f810018", 11263 => x"78010001", 11264 => x"b9601000",
    11265 => x"34030001", 11266 => x"34040000", 11267 => x"38216910",
    11268 => x"fbfffd33", 11269 => x"78020001", 11270 => x"3842808c",
    11271 => x"58410000", 11272 => x"2b9d0004", 11273 => x"2b8b0008",
    11274 => x"379c001c", 11275 => x"c3a00000", 11276 => x"379cffe0",
    11277 => x"5b8b0018", 11278 => x"5b8c0014", 11279 => x"5b8d0010",
    11280 => x"5b8e000c", 11281 => x"5b8f0008", 11282 => x"5b9d0004",
    11283 => x"378d001c", 11284 => x"b8205800", 11285 => x"b9a00800",
    11286 => x"fbffff39", 11287 => x"41620000", 11288 => x"34010045",
    11289 => x"340c0000", 11290 => x"5c41004a", 11291 => x"356e0010",
    11292 => x"b9a01000", 11293 => x"b9c00800", 11294 => x"34030004",
    11295 => x"f8001f83", 11296 => x"b8201000", 11297 => x"5c200043",
    11298 => x"41640009", 11299 => x"34030001", 11300 => x"416d0002",
    11301 => x"41610003", 11302 => x"b8406000", 11303 => x"5c83003d",
    11304 => x"41630014", 11305 => x"34020008", 11306 => x"5c62003a",
    11307 => x"3dad0008", 11308 => x"b9a16800", 11309 => x"35adffe8",
    11310 => x"34010040", 11311 => x"4c2d0002", 11312 => x"340d0040",
    11313 => x"356f000c", 11314 => x"b9e01000", 11315 => x"34030004",
    11316 => x"37810020", 11317 => x"f8001f8e", 11318 => x"35ac0018",
    11319 => x"34010045", 11320 => x"31610000", 11321 => x"15810008",
    11322 => x"3782001c", 11323 => x"31610002", 11324 => x"3401003f",
    11325 => x"31610008", 11326 => x"34010001", 11327 => x"31610009",
    11328 => x"34030004", 11329 => x"31600001", 11330 => x"316c0003",
    11331 => x"31600004", 11332 => x"31600005", 11333 => x"31600006",
    11334 => x"31600007", 11335 => x"3160000a", 11336 => x"3160000b",
    11337 => x"b9e00800", 11338 => x"f8001f79", 11339 => x"34030004",
    11340 => x"37820020", 11341 => x"b9c00800", 11342 => x"f8001f75",
    11343 => x"35ad0005", 11344 => x"01a1001f", 11345 => x"31600014",
    11346 => x"b42d6800", 11347 => x"15a20001", 11348 => x"31600015",
    11349 => x"31600016", 11350 => x"31600017", 11351 => x"35610014",
    11352 => x"fbfffee7", 11353 => x"2021ffff", 11354 => x"00220008",
    11355 => x"31610017", 11356 => x"31620016", 11357 => x"b9600800",
    11358 => x"3402000a", 11359 => x"fbfffee0", 11360 => x"2021ffff",
    11361 => x"00220008", 11362 => x"3161000b", 11363 => x"3162000a",
    11364 => x"b9800800", 11365 => x"2b9d0004", 11366 => x"2b8b0018",
    11367 => x"2b8c0014", 11368 => x"2b8d0010", 11369 => x"2b8e000c",
    11370 => x"2b8f0008", 11371 => x"379c0020", 11372 => x"c3a00000",
    11373 => x"379cffcc", 11374 => x"5b8b0028", 11375 => x"5b8c0024",
    11376 => x"5b8d0020", 11377 => x"5b8e001c", 11378 => x"5b8f0018",
    11379 => x"5b900014", 11380 => x"5b910010", 11381 => x"5b92000c",
    11382 => x"5b930008", 11383 => x"5b9d0004", 11384 => x"b8205800",
    11385 => x"b8406800", 11386 => x"b8606000", 11387 => x"5c600012",
    11388 => x"3562000c", 11389 => x"34030004", 11390 => x"37810030",
    11391 => x"f8001f44", 11392 => x"378c002c", 11393 => x"35620010",
    11394 => x"34030004", 11395 => x"b9800800", 11396 => x"f8001f3f",
    11397 => x"35620014", 11398 => x"34030002", 11399 => x"37810036",
    11400 => x"f8001f3b", 11401 => x"37810034", 11402 => x"35620016",
    11403 => x"34030002", 11404 => x"f8001f37", 11405 => x"35700008",
    11406 => x"b9801000", 11407 => x"34030004", 11408 => x"ba000800",
    11409 => x"f8001f32", 11410 => x"35b1ffec", 11411 => x"356f000c",
    11412 => x"358e0004", 11413 => x"b9c01000", 11414 => x"34030004",
    11415 => x"16320008", 11416 => x"b9e00800", 11417 => x"f8001f2a",
    11418 => x"34010011", 11419 => x"225200ff", 11420 => x"223100ff",
    11421 => x"31610011", 11422 => x"35820008", 11423 => x"34030002",
    11424 => x"31600010", 11425 => x"31720012", 11426 => x"31710013",
    11427 => x"35610014", 11428 => x"f8001f1f", 11429 => x"34030002",
    11430 => x"3582000a", 11431 => x"35610016", 11432 => x"f8001f1b",
    11433 => x"b56d0800", 11434 => x"31720018", 11435 => x"31710019",
    11436 => x"3160001a", 11437 => x"3160001b", 11438 => x"35a2fff9",
    11439 => x"30200000", 11440 => x"0041001f", 11441 => x"35730010",
    11442 => x"b4221000", 11443 => x"14420001", 11444 => x"ba000800",
    11445 => x"fbfffe8a", 11446 => x"2023ffff", 11447 => x"5c600002",
    11448 => x"3803ffff", 11449 => x"00610008", 11450 => x"3163001b",
    11451 => x"3161001a", 11452 => x"34010045", 11453 => x"31610000",
    11454 => x"15a10008", 11455 => x"b9801000", 11456 => x"31610002",
    11457 => x"3401003f", 11458 => x"31610008", 11459 => x"34010011",
    11460 => x"31610009", 11461 => x"31600001", 11462 => x"316d0003",
    11463 => x"31600004", 11464 => x"31600005", 11465 => x"31600006",
    11466 => x"31600007", 11467 => x"3160000a", 11468 => x"3160000b",
    11469 => x"b9e00800", 11470 => x"34030004", 11471 => x"f8001ef4",
    11472 => x"b9c01000", 11473 => x"34030004", 11474 => x"ba600800",
    11475 => x"f8001ef0", 11476 => x"b9600800", 11477 => x"3402000a",
    11478 => x"fbfffe69", 11479 => x"2021ffff", 11480 => x"00220008",
    11481 => x"3161000b", 11482 => x"3162000a", 11483 => x"2b9d0004",
    11484 => x"2b8b0028", 11485 => x"2b8c0024", 11486 => x"2b8d0020",
    11487 => x"2b8e001c", 11488 => x"2b8f0018", 11489 => x"2b900014",
    11490 => x"2b910010", 11491 => x"2b92000c", 11492 => x"2b930008",
    11493 => x"379c0034", 11494 => x"c3a00000", 11495 => x"379cffe4",
    11496 => x"5b8b0010", 11497 => x"5b8c000c", 11498 => x"5b8d0008",
    11499 => x"5b9d0004", 11500 => x"b8405800", 11501 => x"b8206800",
    11502 => x"34020001", 11503 => x"34010006", 11504 => x"3162001c",
    11505 => x"3162001d", 11506 => x"3161001e", 11507 => x"3160001f",
    11508 => x"35610020", 11509 => x"b8606000", 11510 => x"f8000601",
    11511 => x"41620024", 11512 => x"41610020", 11513 => x"34030002",
    11514 => x"98410800", 11515 => x"31610020", 11516 => x"41620025",
    11517 => x"41610021", 11518 => x"316c0025", 11519 => x"98410800",
    11520 => x"31610021", 11521 => x"41610022", 11522 => x"15820008",
    11523 => x"98410800", 11524 => x"31610022", 11525 => x"41610023",
    11526 => x"31620024", 11527 => x"34020000", 11528 => x"982c0800",
    11529 => x"31610023", 11530 => x"35610026", 11531 => x"f8001f36",
    11532 => x"35610028", 11533 => x"34020000", 11534 => x"34030004",
    11535 => x"f8001f32", 11536 => x"3561002c", 11537 => x"34020000",
    11538 => x"34030004", 11539 => x"f8001f2e", 11540 => x"35610030",
    11541 => x"34020000", 11542 => x"34030004", 11543 => x"f8001f2a",
    11544 => x"35610034", 11545 => x"34020000", 11546 => x"34030004",
    11547 => x"f8001f26", 11548 => x"356c0038", 11549 => x"34020000",
    11550 => x"34030010", 11551 => x"b9800800", 11552 => x"f8001f21",
    11553 => x"b9800800", 11554 => x"f80005d5", 11555 => x"35610048",
    11556 => x"34020000", 11557 => x"34030040", 11558 => x"f8001f1b",
    11559 => x"35610088", 11560 => x"34020000", 11561 => x"34030080",
    11562 => x"f8001f17", 11563 => x"35610108", 11564 => x"34020000",
    11565 => x"34030040", 11566 => x"f8001f13", 11567 => x"378c0014",
    11568 => x"b9800800", 11569 => x"34020000", 11570 => x"34030004",
    11571 => x"f8001f0e", 11572 => x"37810018", 11573 => x"340200ff",
    11574 => x"34030004", 11575 => x"f8001f0a", 11576 => x"34010044",
    11577 => x"0f81001c", 11578 => x"34010043", 11579 => x"0f81001e",
    11580 => x"b9801800", 11581 => x"b9600800", 11582 => x"34020148",
    11583 => x"fbffff2e", 11584 => x"b9a00800", 11585 => x"340200ff",
    11586 => x"34030006", 11587 => x"f8001efe", 11588 => x"34010148",
    11589 => x"2b9d0004", 11590 => x"2b8b0010", 11591 => x"2b8c000c",
    11592 => x"2b8d0008", 11593 => x"379c001c", 11594 => x"c3a00000",
    11595 => x"379cffe0", 11596 => x"5b8b0014", 11597 => x"5b8c0010",
    11598 => x"5b8d000c", 11599 => x"5b8e0008", 11600 => x"5b9d0004",
    11601 => x"378d0018", 11602 => x"b8205800", 11603 => x"b9a00800",
    11604 => x"b8407000", 11605 => x"f80005a2", 11606 => x"34010148",
    11607 => x"340c0000", 11608 => x"5dc1001b", 11609 => x"41610014",
    11610 => x"5c200019", 11611 => x"41620015", 11612 => x"34010043",
    11613 => x"5c410016", 11614 => x"35610038", 11615 => x"b9a01000",
    11616 => x"34030006", 11617 => x"f8001e41", 11618 => x"5c200011",
    11619 => x"78010001", 11620 => x"34020001", 11621 => x"38217d90",
    11622 => x"58220000", 11623 => x"3561002c", 11624 => x"fbfffdf0",
    11625 => x"37810020", 11626 => x"fbfffde5", 11627 => x"43820020",
    11628 => x"43830021", 11629 => x"43840022", 11630 => x"43850023",
    11631 => x"78010001", 11632 => x"3821559c", 11633 => x"f800047e",
    11634 => x"340c0001", 11635 => x"b9800800", 11636 => x"2b9d0004",
    11637 => x"2b8b0014", 11638 => x"2b8c0010", 11639 => x"2b8d000c",
    11640 => x"2b8e0008", 11641 => x"379c0020", 11642 => x"c3a00000",
    11643 => x"379cfffc", 11644 => x"5b8b0004", 11645 => x"78040001",
    11646 => x"38845e2c", 11647 => x"3442ffff", 11648 => x"348a001c",
    11649 => x"34030000", 11650 => x"340900fd", 11651 => x"340800f9",
    11652 => x"340700ff", 11653 => x"3406ffa2", 11654 => x"e0000011",
    11655 => x"40850000", 11656 => x"5ca90004", 11657 => x"b4232800",
    11658 => x"30a60000", 11659 => x"e000000a", 11660 => x"5ca80005",
    11661 => x"b4232800", 11662 => x"40a50000", 11663 => x"b4651800",
    11664 => x"e0000005", 11665 => x"5ca70004", 11666 => x"b4232800",
    11667 => x"c8435800", 11668 => x"30ab0000", 11669 => x"34630001",
    11670 => x"34840001", 11671 => x"5c8afff0", 11672 => x"2b8b0004",
    11673 => x"379c0004", 11674 => x"c3a00000", 11675 => x"379cfff8",
    11676 => x"5b8b0008", 11677 => x"5b9d0004", 11678 => x"40230006",
    11679 => x"34040020", 11680 => x"4c830002", 11681 => x"34030020",
    11682 => x"206b00ff", 11683 => x"b42b1800", 11684 => x"3404ffa2",
    11685 => x"30640007", 11686 => x"4063000a", 11687 => x"34040004",
    11688 => x"4c830002", 11689 => x"34030004", 11690 => x"b5635800",
    11691 => x"216b00ff", 11692 => x"b42b1800", 11693 => x"3062000d",
    11694 => x"34020001", 11695 => x"30620010", 11696 => x"40620016",
    11697 => x"34030028", 11698 => x"4c620002", 11699 => x"34020028",
    11700 => x"b5621000", 11701 => x"204200ff", 11702 => x"b4221800",
    11703 => x"34420019", 11704 => x"34040005", 11705 => x"204b00ff",
    11706 => x"30640017", 11707 => x"30600018", 11708 => x"b9601000",
    11709 => x"fbffffbe", 11710 => x"b9600800", 11711 => x"2b9d0004",
    11712 => x"2b8b0008", 11713 => x"379c0008", 11714 => x"c3a00000",
    11715 => x"379cfefc", 11716 => x"5b8b0028", 11717 => x"5b8c0024",
    11718 => x"5b8d0020", 11719 => x"5b8e001c", 11720 => x"5b8f0018",
    11721 => x"5b900014", 11722 => x"5b910010", 11723 => x"5b92000c",
    11724 => x"5b930008", 11725 => x"5b9d0004", 11726 => x"78010001",
    11727 => x"38218110", 11728 => x"28210000", 11729 => x"378b002c",
    11730 => x"378200f4", 11731 => x"b9601800", 11732 => x"340400c8",
    11733 => x"34050000", 11734 => x"fbfffc04", 11735 => x"34020038",
    11736 => x"340c0000", 11737 => x"504100a6", 11738 => x"b9600800",
    11739 => x"fbfffda6", 11740 => x"5c2000a3", 11741 => x"78010001",
    11742 => x"78020001", 11743 => x"38219298", 11744 => x"38425e2c",
    11745 => x"78030001", 11746 => x"40250000", 11747 => x"344e001c",
    11748 => x"b9600800", 11749 => x"34040000", 11750 => x"340d0006",
    11751 => x"38635e10", 11752 => x"340b00a0", 11753 => x"340a00a1",
    11754 => x"340900a3", 11755 => x"34080001", 11756 => x"e0000028",
    11757 => x"40460000", 11758 => x"34c70007", 11759 => x"20e700ff",
    11760 => x"54ed0014", 11761 => x"3ce70002", 11762 => x"b4673800",
    11763 => x"28e60000", 11764 => x"c0c00000", 11765 => x"b4813000",
    11766 => x"40c6001c", 11767 => x"b4862000", 11768 => x"e000001a",
    11769 => x"b4812800", 11770 => x"40a5001c", 11771 => x"51050017",
    11772 => x"e000000b", 11773 => x"b4813000", 11774 => x"40c6001c",
    11775 => x"44cb000e", 11776 => x"44ca000f", 11777 => x"44c90010",
    11778 => x"5d800010", 11779 => x"e0000004", 11780 => x"b4813800",
    11781 => x"40e7001c", 11782 => x"44e6000c", 11783 => x"78010001",
    11784 => x"38219298", 11785 => x"30250000", 11786 => x"34020005",
    11787 => x"37810048", 11788 => x"e000005b", 11789 => x"340c0002",
    11790 => x"e0000004", 11791 => x"340c0004", 11792 => x"e0000002",
    11793 => x"340c0001", 11794 => x"34840001", 11795 => x"34420001",
    11796 => x"5c4effd9", 11797 => x"78010001", 11798 => x"38219298",
    11799 => x"30250000", 11800 => x"37810048", 11801 => x"b4246800",
    11802 => x"780b0001", 11803 => x"34840001", 11804 => x"b4247800",
    11805 => x"396b6964", 11806 => x"21930003", 11807 => x"21900004",
    11808 => x"39920008", 11809 => x"e000003f", 11810 => x"41b10000",
    11811 => x"46600002", 11812 => x"5431003b", 11813 => x"222200ff",
    11814 => x"50220002", 11815 => x"b8208800", 11816 => x"29610000",
    11817 => x"223100ff", 11818 => x"b9e01000", 11819 => x"ba201800",
    11820 => x"f8001d76", 11821 => x"3c250018", 11822 => x"b9807000",
    11823 => x"14a50018", 11824 => x"4600000a", 11825 => x"48a00007",
    11826 => x"4163000c", 11827 => x"41a10000", 11828 => x"64a20000",
    11829 => x"f0610800", 11830 => x"a0410800", 11831 => x"44200003",
    11832 => x"4171000c", 11833 => x"ba407000", 11834 => x"4163000c",
    11835 => x"64a10000", 11836 => x"e4711000", 11837 => x"a0411000",
    11838 => x"5c400003", 11839 => x"21c10008", 11840 => x"4422001e",
    11841 => x"5e000003", 11842 => x"21c10008", 11843 => x"44300004",
    11844 => x"29620000", 11845 => x"b9e00800", 11846 => x"f8001d7d",
    11847 => x"29650004", 11848 => x"29630008", 11849 => x"b9a00800",
    11850 => x"ba201000", 11851 => x"b9c02000", 11852 => x"d8a00000",
    11853 => x"4c01000c", 11854 => x"5e000003", 11855 => x"21ce0008",
    11856 => x"45d00005", 11857 => x"41a30000", 11858 => x"4162000c",
    11859 => x"b4621000", 11860 => x"31a20000", 11861 => x"4164000c",
    11862 => x"b5e47800", 11863 => x"b5e17800", 11864 => x"e000000a",
    11865 => x"44200006", 11866 => x"c8011000", 11867 => x"204200ff",
    11868 => x"37810048", 11869 => x"e000000a", 11870 => x"48a10007",
    11871 => x"356b0010", 11872 => x"4161000c", 11873 => x"5c20ffc1",
    11874 => x"45600003", 11875 => x"4161000c", 11876 => x"5c200006",
    11877 => x"37810048", 11878 => x"34020002", 11879 => x"fbffff34",
    11880 => x"b8205800", 11881 => x"e0000007", 11882 => x"37810048",
    11883 => x"c9e15800", 11884 => x"b9601000", 11885 => x"fbffff0e",
    11886 => x"340c0000", 11887 => x"480b0010", 11888 => x"378c002c",
    11889 => x"356b001c", 11890 => x"b9800800", 11891 => x"b9601000",
    11892 => x"34030000", 11893 => x"fbfffdf8", 11894 => x"78050001",
    11895 => x"38a58110", 11896 => x"28a10000", 11897 => x"b9801800",
    11898 => x"378200f4", 11899 => x"b9602000", 11900 => x"34050000",
    11901 => x"fbfffbcf", 11902 => x"340c0001", 11903 => x"b9800800",
    11904 => x"2b9d0004", 11905 => x"2b8b0028", 11906 => x"2b8c0024",
    11907 => x"2b8d0020", 11908 => x"2b8e001c", 11909 => x"2b8f0018",
    11910 => x"2b900014", 11911 => x"2b910010", 11912 => x"2b92000c",
    11913 => x"2b930008", 11914 => x"379c0104", 11915 => x"c3a00000",
    11916 => x"379cffec", 11917 => x"5b8b0010", 11918 => x"5b8c000c",
    11919 => x"5b8d0008", 11920 => x"5b9d0004", 11921 => x"b8403000",
    11922 => x"40c50011", 11923 => x"40220000", 11924 => x"b8606000",
    11925 => x"402b0001", 11926 => x"3404fffd", 11927 => x"5ca2001e",
    11928 => x"34220002", 11929 => x"34010004", 11930 => x"44a10013",
    11931 => x"34010042", 11932 => x"44a10004", 11933 => x"34010002",
    11934 => x"34040000", 11935 => x"5ca10016", 11936 => x"340d0004",
    11937 => x"3404fffd", 11938 => x"556d0013", 11939 => x"37810014",
    11940 => x"b9601800", 11941 => x"5b800014", 11942 => x"f8001d1d",
    11943 => x"2b810014", 11944 => x"c9ab6800", 11945 => x"3dad0003",
    11946 => x"802d6800", 11947 => x"598d0000", 11948 => x"e0000008",
    11949 => x"40c10013", 11950 => x"55610007", 11951 => x"b8600800",
    11952 => x"b58b6000", 11953 => x"b9601800", 11954 => x"f8001d11",
    11955 => x"31800000", 11956 => x"35640002", 11957 => x"b8800800",
    11958 => x"2b9d0004", 11959 => x"2b8b0010", 11960 => x"2b8c000c",
    11961 => x"2b8d0008", 11962 => x"379c0014", 11963 => x"c3a00000",
    11964 => x"379cfffc", 11965 => x"5b9d0004", 11966 => x"40430012",
    11967 => x"2844000c", 11968 => x"b4831800", 11969 => x"fbffffcb",
    11970 => x"2b9d0004", 11971 => x"379c0004", 11972 => x"c3a00000",
    11973 => x"379cffcc", 11974 => x"5b8b0020", 11975 => x"5b8c001c",
    11976 => x"5b8d0018", 11977 => x"5b8e0014", 11978 => x"5b8f0010",
    11979 => x"5b90000c", 11980 => x"5b910008", 11981 => x"5b9d0004",
    11982 => x"402e0000", 11983 => x"204200ff", 11984 => x"208400ff",
    11985 => x"344c0001", 11986 => x"c9c27000", 11987 => x"20820001",
    11988 => x"b8207800", 11989 => x"b42c6000", 11990 => x"3401fffc",
    11991 => x"5c400068", 11992 => x"208d0004", 11993 => x"7dad0000",
    11994 => x"20900008", 11995 => x"7e100000", 11996 => x"b8605800",
    11997 => x"21b100ff", 11998 => x"e0000023", 11999 => x"b9c01800",
    12000 => x"4c2e0002", 12001 => x"b8201800", 12002 => x"29610000",
    12003 => x"b9801000", 12004 => x"206300ff", 12005 => x"f8001cbd",
    12006 => x"5e00000a", 12007 => x"b0200800", 12008 => x"64220000",
    12009 => x"a0511800", 12010 => x"44700003", 12011 => x"41630010",
    12012 => x"4c6e0004", 12013 => x"68210000", 12014 => x"a2210800",
    12015 => x"4420000b", 12016 => x"29620000", 12017 => x"41630010",
    12018 => x"b9800800", 12019 => x"340e0000", 12020 => x"f8001ccf",
    12021 => x"41610010", 12022 => x"34020001", 12023 => x"b5810800",
    12024 => x"30220000", 12025 => x"e000000d", 12026 => x"44410006",
    12027 => x"41610010", 12028 => x"34210001", 12029 => x"45c10006",
    12030 => x"45a00002", 12031 => x"49c10006", 12032 => x"356b0014",
    12033 => x"41610010", 12034 => x"5c20ffdd", 12035 => x"b9a07000",
    12036 => x"e0000002", 12037 => x"340e0001", 12038 => x"41620010",
    12039 => x"34010000", 12040 => x"44400037", 12041 => x"41610011",
    12042 => x"33820034", 12043 => x"5b8c0024", 12044 => x"33810035",
    12045 => x"2961000c", 12046 => x"5b810030", 12047 => x"45c00004",
    12048 => x"41810001", 12049 => x"34210001", 12050 => x"31810001",
    12051 => x"41610010", 12052 => x"29630004", 12053 => x"37910024",
    12054 => x"34210001", 12055 => x"b5810800", 12056 => x"ba201000",
    12057 => x"d8600000", 12058 => x"64230000", 12059 => x"a06e7000",
    12060 => x"45c00019", 12061 => x"356b0014", 12062 => x"41630010",
    12063 => x"34010000", 12064 => x"4460001f", 12065 => x"29620000",
    12066 => x"b9800800", 12067 => x"f8001ca0", 12068 => x"41610010",
    12069 => x"34020001", 12070 => x"b5810800", 12071 => x"30220000",
    12072 => x"41620011", 12073 => x"41610010", 12074 => x"29630004",
    12075 => x"33820035", 12076 => x"2962000c", 12077 => x"33810034",
    12078 => x"34210001", 12079 => x"5b820030", 12080 => x"b5810800",
    12081 => x"ba201000", 12082 => x"d8600000", 12083 => x"5c200003",
    12084 => x"e000000b", 12085 => x"5c6e0009", 12086 => x"48010009",
    12087 => x"41620010", 12088 => x"ba0d6800", 12089 => x"34420001",
    12090 => x"b4220800", 12091 => x"45a00004", 12092 => x"31e20000",
    12093 => x"e0000002", 12094 => x"34010000", 12095 => x"2b9d0004",
    12096 => x"2b8b0020", 12097 => x"2b8c001c", 12098 => x"2b8d0018",
    12099 => x"2b8e0014", 12100 => x"2b8f0010", 12101 => x"2b90000c",
    12102 => x"2b910008", 12103 => x"379c0034", 12104 => x"c3a00000",
    12105 => x"379cffd0", 12106 => x"5b8b0030", 12107 => x"5b8c002c",
    12108 => x"5b8d0028", 12109 => x"5b8e0024", 12110 => x"5b8f0020",
    12111 => x"5b90001c", 12112 => x"5b910018", 12113 => x"5b920014",
    12114 => x"5b930010", 12115 => x"5b94000c", 12116 => x"5b950008",
    12117 => x"5b9d0004", 12118 => x"208400ff", 12119 => x"40310000",
    12120 => x"204200ff", 12121 => x"008d0003", 12122 => x"344e0001",
    12123 => x"208f0004", 12124 => x"b8208000", 12125 => x"ca228800",
    12126 => x"b42e7000", 12127 => x"21ad0001", 12128 => x"b8605800",
    12129 => x"340c0000", 12130 => x"20950003", 12131 => x"20940001",
    12132 => x"7df30000", 12133 => x"e0000034", 12134 => x"b8a09000",
    12135 => x"5da00005", 12136 => x"ba209000", 12137 => x"4cb10002",
    12138 => x"b8a09000", 12139 => x"225200ff", 12140 => x"46a00002",
    12141 => x"5e25002b", 12142 => x"5da0000c", 12143 => x"29610000",
    12144 => x"b9c01000", 12145 => x"ba401800", 12146 => x"f8001c30",
    12147 => x"3c2c0018", 12148 => x"158c0018", 12149 => x"5d8d0006",
    12150 => x"45ec0009", 12151 => x"41610010", 12152 => x"5c320007",
    12153 => x"e000001f", 12154 => x"45800005", 12155 => x"69810000",
    12156 => x"a0331000", 12157 => x"5c400002", 12158 => x"45a20019",
    12159 => x"45e00007", 12160 => x"29620000", 12161 => x"41630010",
    12162 => x"b9c00800", 12163 => x"f8001c40", 12164 => x"41610010",
    12165 => x"32010000", 12166 => x"46800008", 12167 => x"29630008",
    12168 => x"44600014", 12169 => x"41610010", 12170 => x"b9601000",
    12171 => x"b5c10800", 12172 => x"d8600000", 12173 => x"48010012",
    12174 => x"41610010", 12175 => x"29630004", 12176 => x"b9601000",
    12177 => x"b5c10800", 12178 => x"d8600000", 12179 => x"44200005",
    12180 => x"41620010", 12181 => x"b4220800", 12182 => x"e0000009",
    12183 => x"5c2d0007", 12184 => x"356b0014", 12185 => x"41650010",
    12186 => x"5ca0ffcc", 12187 => x"e0000003", 12188 => x"3401fffc",
    12189 => x"e0000002", 12190 => x"34010000", 12191 => x"2b9d0004",
    12192 => x"2b8b0030", 12193 => x"2b8c002c", 12194 => x"2b8d0028",
    12195 => x"2b8e0024", 12196 => x"2b8f0020", 12197 => x"2b90001c",
    12198 => x"2b910018", 12199 => x"2b920014", 12200 => x"2b930010",
    12201 => x"2b94000c", 12202 => x"2b950008", 12203 => x"379c0030",
    12204 => x"c3a00000", 12205 => x"379cffe4", 12206 => x"5b8b0010",
    12207 => x"5b8c000c", 12208 => x"5b8d0008", 12209 => x"5b9d0004",
    12210 => x"b8206000", 12211 => x"342d0002", 12212 => x"30220000",
    12213 => x"34010043", 12214 => x"b8605800", 12215 => x"54410008",
    12216 => x"34010041", 12217 => x"50410009", 12218 => x"34010002",
    12219 => x"44410007", 12220 => x"34010004", 12221 => x"5c410029",
    12222 => x"e000001c", 12223 => x"34010046", 12224 => x"5c410026",
    12225 => x"e0000009", 12226 => x"29610000", 12227 => x"3782001c",
    12228 => x"34030004", 12229 => x"5b81001c", 12230 => x"b9a00800",
    12231 => x"f8001bfc", 12232 => x"34010004", 12233 => x"e000000f",
    12234 => x"78010001", 12235 => x"38219298", 12236 => x"40210000",
    12237 => x"34020000", 12238 => x"44200019", 12239 => x"28610000",
    12240 => x"37820014", 12241 => x"5b810014", 12242 => x"28610004",
    12243 => x"34030008", 12244 => x"5b810018", 12245 => x"b9a00800",
    12246 => x"f8001bed", 12247 => x"34010008", 12248 => x"31810001",
    12249 => x"e000000a", 12250 => x"b8600800", 12251 => x"3402001f",
    12252 => x"f8001dca", 12253 => x"202300ff", 12254 => x"31830001",
    12255 => x"b9a00800", 12256 => x"b9601000", 12257 => x"34630001",
    12258 => x"f8001be1", 12259 => x"41820001", 12260 => x"34420002",
    12261 => x"e0000002", 12262 => x"34020000", 12263 => x"b8400800",
    12264 => x"2b9d0004", 12265 => x"2b8b0010", 12266 => x"2b8c000c",
    12267 => x"2b8d0008", 12268 => x"379c001c", 12269 => x"c3a00000",
    12270 => x"379cff98", 12271 => x"5b8b0034", 12272 => x"5b8c0030",
    12273 => x"5b8d002c", 12274 => x"5b8e0028", 12275 => x"5b8f0024",
    12276 => x"5b900020", 12277 => x"5b91001c", 12278 => x"5b920018",
    12279 => x"5b930014", 12280 => x"5b940010", 12281 => x"5b95000c",
    12282 => x"5b960008", 12283 => x"5b9d0004", 12284 => x"b8208000",
    12285 => x"28410000", 12286 => x"b8407000", 12287 => x"340d0000",
    12288 => x"40360001", 12289 => x"402c0000", 12290 => x"340b0001",
    12291 => x"378f0038", 12292 => x"3415ffff", 12293 => x"34140002",
    12294 => x"34130003", 12295 => x"34120004", 12296 => x"34110005",
    12297 => x"21a300ff", 12298 => x"b9e00800", 12299 => x"34020000",
    12300 => x"f8000c39", 12301 => x"b8201800", 12302 => x"4420001c",
    12303 => x"4435001b", 12304 => x"5ecb000d", 12305 => x"5d940009",
    12306 => x"378b0058", 12307 => x"34030010", 12308 => x"b9600800",
    12309 => x"b9e01000", 12310 => x"f8001bad", 12311 => x"b9601800",
    12312 => x"33800068", 12313 => x"e000000d", 12314 => x"45930007",
    12315 => x"45920008", 12316 => x"45910009", 12317 => x"356b0001",
    12318 => x"35ad0001", 12319 => x"4c6bffea", 12320 => x"e000000a",
    12321 => x"3783004c", 12322 => x"e0000004", 12323 => x"37830050",
    12324 => x"e0000002", 12325 => x"37830048", 12326 => x"41c20011",
    12327 => x"ba000800", 12328 => x"fbffff85", 12329 => x"e0000002",
    12330 => x"34010000", 12331 => x"2b9d0004", 12332 => x"2b8b0034",
    12333 => x"2b8c0030", 12334 => x"2b8d002c", 12335 => x"2b8e0028",
    12336 => x"2b8f0024", 12337 => x"2b900020", 12338 => x"2b91001c",
    12339 => x"2b920018", 12340 => x"2b930014", 12341 => x"2b940010",
    12342 => x"2b95000c", 12343 => x"2b960008", 12344 => x"379c0068",
    12345 => x"c3a00000", 12346 => x"379cffe8", 12347 => x"5b8b0010",
    12348 => x"5b8c000c", 12349 => x"5b8d0008", 12350 => x"5b9d0004",
    12351 => x"b8405800", 12352 => x"2842000c", 12353 => x"34030001",
    12354 => x"b8206800", 12355 => x"44430019", 12356 => x"34030002",
    12357 => x"5c43002e", 12358 => x"78020001", 12359 => x"38428114",
    12360 => x"28430000", 12361 => x"286400b4", 12362 => x"286500b0",
    12363 => x"c8042000", 12364 => x"7c820000", 12365 => x"c8052800",
    12366 => x"c8a22800", 12367 => x"3c820001", 12368 => x"3ca50001",
    12369 => x"f4822000", 12370 => x"b4852000", 12371 => x"286500a0",
    12372 => x"286300a4", 12373 => x"b4852000", 12374 => x"b4431800",
    12375 => x"f4431000", 12376 => x"5b830018", 12377 => x"b4441000",
    12378 => x"5b820014", 12379 => x"e0000014", 12380 => x"78020001",
    12381 => x"38428114", 12382 => x"284c0000", 12383 => x"78050001",
    12384 => x"38a55a2c", 12385 => x"298200fc", 12386 => x"28a40000",
    12387 => x"34030000", 12388 => x"1441001f", 12389 => x"f8001a89",
    12390 => x"29830100", 12391 => x"1464001f", 12392 => x"b4431800",
    12393 => x"f4431000", 12394 => x"b4242000", 12395 => x"b4442000",
    12396 => x"5b840014", 12397 => x"5b830018", 12398 => x"b9a00800",
    12399 => x"41620011", 12400 => x"37830014", 12401 => x"fbffff3c",
    12402 => x"e0000002", 12403 => x"3401ffff", 12404 => x"2b9d0004",
    12405 => x"2b8b0010", 12406 => x"2b8c000c", 12407 => x"2b8d0008",
    12408 => x"379c0018", 12409 => x"c3a00000", 12410 => x"379cfff8",
    12411 => x"5b9d0004", 12412 => x"2843000c", 12413 => x"40450011",
    12414 => x"40420012", 12415 => x"28630000", 12416 => x"b4621000",
    12417 => x"28440000", 12418 => x"28430004", 12419 => x"4880000e",
    12420 => x"5c800005", 12421 => x"78060001", 12422 => x"38c65a44",
    12423 => x"28c20000", 12424 => x"54620009", 12425 => x"3402ffff",
    12426 => x"4844000b", 12427 => x"5c82000b", 12428 => x"78040001",
    12429 => x"38845a48", 12430 => x"28820000", 12431 => x"54430006",
    12432 => x"e0000006", 12433 => x"78060001", 12434 => x"38c65a68",
    12435 => x"28c30000", 12436 => x"e0000002", 12437 => x"78038000",
    12438 => x"5b830008", 12439 => x"b8a01000", 12440 => x"37830008",
    12441 => x"fbffff14", 12442 => x"2b9d0004", 12443 => x"379c0008",
    12444 => x"c3a00000", 12445 => x"379cfffc", 12446 => x"5b9d0004",
    12447 => x"2844000c", 12448 => x"40430012", 12449 => x"40420011",
    12450 => x"28840000", 12451 => x"b4831800", 12452 => x"fbffff09",
    12453 => x"2b9d0004", 12454 => x"379c0004", 12455 => x"c3a00000",
    12456 => x"379cfffc", 12457 => x"5b9d0004", 12458 => x"2844000c",
    12459 => x"40430012", 12460 => x"40420011", 12461 => x"b4831800",
    12462 => x"fbfffeff", 12463 => x"2b9d0004", 12464 => x"379c0004",
    12465 => x"c3a00000", 12466 => x"379cfff0", 12467 => x"5b8b000c",
    12468 => x"5b8c0008", 12469 => x"5b9d0004", 12470 => x"b8405800",
    12471 => x"2842000c", 12472 => x"b8206000", 12473 => x"34010001",
    12474 => x"5c41000a", 12475 => x"34010000", 12476 => x"f8000286",
    12477 => x"34220001", 12478 => x"5b820010", 12479 => x"41620011",
    12480 => x"b9800800", 12481 => x"37830010", 12482 => x"fbfffeeb",
    12483 => x"e0000002", 12484 => x"3401ffff", 12485 => x"2b9d0004",
    12486 => x"2b8b000c", 12487 => x"2b8c0008", 12488 => x"379c0010",
    12489 => x"c3a00000", 12490 => x"379cfff4", 12491 => x"5b8b000c",
    12492 => x"5b8c0008", 12493 => x"5b9d0004", 12494 => x"284b000c",
    12495 => x"b9601800", 12496 => x"fbfffdbc", 12497 => x"b8206000",
    12498 => x"4c01000a", 12499 => x"29620000", 12500 => x"34010001",
    12501 => x"5c410005", 12502 => x"fbffd2c3", 12503 => x"fbffd29c",
    12504 => x"34010064", 12505 => x"e0000002", 12506 => x"340100c8",
    12507 => x"59610000", 12508 => x"b9800800", 12509 => x"2b9d0004",
    12510 => x"2b8b000c", 12511 => x"2b8c0008", 12512 => x"379c000c",
    12513 => x"c3a00000", 12514 => x"379cfff0", 12515 => x"5b8b0010",
    12516 => x"5b8c000c", 12517 => x"5b8d0008", 12518 => x"5b9d0004",
    12519 => x"284b000c", 12520 => x"b9601800", 12521 => x"fbfffda3",
    12522 => x"b8206800", 12523 => x"4c010050", 12524 => x"29620000",
    12525 => x"34010002", 12526 => x"4441001e", 12527 => x"48410004",
    12528 => x"34010001", 12529 => x"5c410048", 12530 => x"e0000020",
    12531 => x"34010003", 12532 => x"44410004", 12533 => x"34010032",
    12534 => x"5c410043", 12535 => x"e000003d", 12536 => x"78020001",
    12537 => x"38428118", 12538 => x"28410014", 12539 => x"78030001",
    12540 => x"38638ec8", 12541 => x"58610000", 12542 => x"28410018",
    12543 => x"78030001", 12544 => x"38638ecc", 12545 => x"58610000",
    12546 => x"28410010", 12547 => x"78030001", 12548 => x"38636ffc",
    12549 => x"58610000", 12550 => x"78010001", 12551 => x"382155c4",
    12552 => x"f80000e7", 12553 => x"fbffd290", 12554 => x"fbffd269",
    12555 => x"e000002c", 12556 => x"78010001", 12557 => x"78020001",
    12558 => x"38218118", 12559 => x"38428f34", 12560 => x"34030010",
    12561 => x"f8001ab2", 12562 => x"780c0001", 12563 => x"398c8118",
    12564 => x"41810000", 12565 => x"5c200003", 12566 => x"340100cb",
    12567 => x"e0000023", 12568 => x"34020010", 12569 => x"b9800800",
    12570 => x"f8001c8c", 12571 => x"b8201000", 12572 => x"3403000f",
    12573 => x"34010020", 12574 => x"e0000004", 12575 => x"b44c2000",
    12576 => x"30810000", 12577 => x"34420001", 12578 => x"4c62fffd",
    12579 => x"34020001", 12580 => x"b9800800", 12581 => x"34030000",
    12582 => x"f8000b1f", 12583 => x"b8201000", 12584 => x"3401fffe",
    12585 => x"5c410003", 12586 => x"340100ca", 12587 => x"e000000f",
    12588 => x"3401ffff", 12589 => x"5c410003", 12590 => x"340100c9",
    12591 => x"e000000b", 12592 => x"f80006da", 12593 => x"44200006",
    12594 => x"34010065", 12595 => x"e0000007", 12596 => x"f8000af8",
    12597 => x"3402ffff", 12598 => x"44220003", 12599 => x"34010064",
    12600 => x"e0000002", 12601 => x"340100c8", 12602 => x"59610000",
    12603 => x"b9a00800", 12604 => x"2b9d0004", 12605 => x"2b8b0010",
    12606 => x"2b8c000c", 12607 => x"2b8d0008", 12608 => x"379c0010",
    12609 => x"c3a00000", 12610 => x"379cffc8", 12611 => x"5b8b0024",
    12612 => x"5b8c0020", 12613 => x"5b8d001c", 12614 => x"5b8e0018",
    12615 => x"5b8f0014", 12616 => x"5b900010", 12617 => x"5b91000c",
    12618 => x"5b920008", 12619 => x"5b9d0004", 12620 => x"b8207800",
    12621 => x"28410000", 12622 => x"b8406800", 12623 => x"340c0001",
    12624 => x"40320001", 12625 => x"402e0000", 12626 => x"34010000",
    12627 => x"f8000913", 12628 => x"b8202000", 12629 => x"34110002",
    12630 => x"34100003", 12631 => x"e0000025", 12632 => x"5e4c0020",
    12633 => x"288b0004", 12634 => x"5dd10007", 12635 => x"28830000",
    12636 => x"78020001", 12637 => x"37810028", 12638 => x"38424aa4",
    12639 => x"f8000082", 12640 => x"e000001f", 12641 => x"5dd00017",
    12642 => x"78018000", 12643 => x"5d610006", 12644 => x"78020001",
    12645 => x"37810028", 12646 => x"384255f0", 12647 => x"f800007a",
    12648 => x"e0000017", 12649 => x"4d600006", 12650 => x"78020001",
    12651 => x"37810028", 12652 => x"3842469c", 12653 => x"c80b5800",
    12654 => x"f8000073", 12655 => x"2164ffff", 12656 => x"08842710",
    12657 => x"78020001", 12658 => x"15630010", 12659 => x"00840010",
    12660 => x"37810028", 12661 => x"384255f8", 12662 => x"f800006b",
    12663 => x"e0000008", 12664 => x"b8800800", 12665 => x"f80008ed",
    12666 => x"b8202000", 12667 => x"358c0001", 12668 => x"5c80ffdc",
    12669 => x"34010000", 12670 => x"e0000005", 12671 => x"41a20011",
    12672 => x"b9e00800", 12673 => x"37830028", 12674 => x"fbfffe2b",
    12675 => x"2b9d0004", 12676 => x"2b8b0024", 12677 => x"2b8c0020",
    12678 => x"2b8d001c", 12679 => x"2b8e0018", 12680 => x"2b8f0014",
    12681 => x"2b900010", 12682 => x"2b91000c", 12683 => x"2b920008",
    12684 => x"379c0038", 12685 => x"c3a00000", 12686 => x"379cffe4",
    12687 => x"5b8b0010", 12688 => x"5b8c000c", 12689 => x"5b8d0008",
    12690 => x"5b9d0004", 12691 => x"284d000c", 12692 => x"b8206000",
    12693 => x"b8405800", 12694 => x"21a10002", 12695 => x"44200009",
    12696 => x"f8000617", 12697 => x"3402000a", 12698 => x"f80019c8",
    12699 => x"5b81001c", 12700 => x"41620011", 12701 => x"b9800800",
    12702 => x"3783001c", 12703 => x"e0000013", 12704 => x"21a20004",
    12705 => x"44410004", 12706 => x"37810014", 12707 => x"34020000",
    12708 => x"f80009a7", 12709 => x"21ad0001", 12710 => x"45a00009",
    12711 => x"2b820018", 12712 => x"2b810014", 12713 => x"34030002",
    12714 => x"fbfff565", 12715 => x"b8201800", 12716 => x"41620011",
    12717 => x"b9800800", 12718 => x"e0000004", 12719 => x"41620011",
    12720 => x"b9800800", 12721 => x"37830014", 12722 => x"fbfffdfb",
    12723 => x"2b9d0004", 12724 => x"2b8b0010", 12725 => x"2b8c000c",
    12726 => x"2b8d0008", 12727 => x"379c001c", 12728 => x"c3a00000",
    12729 => x"379cfffc", 12730 => x"5b9d0004", 12731 => x"78010001",
    12732 => x"34020000", 12733 => x"34030000", 12734 => x"340400a1",
    12735 => x"382169f4", 12736 => x"fbfff777", 12737 => x"78020001",
    12738 => x"38428110", 12739 => x"58410000", 12740 => x"78010001",
    12741 => x"38216178", 12742 => x"28210014", 12743 => x"78020001",
    12744 => x"38428114", 12745 => x"58410000", 12746 => x"2b9d0004",
    12747 => x"379c0004", 12748 => x"c3a00000", 12749 => x"379cfff4",
    12750 => x"5b8b000c", 12751 => x"5b8c0008", 12752 => x"5b9d0004",
    12753 => x"780b0001", 12754 => x"b8202000", 12755 => x"396b8240",
    12756 => x"b8401800", 12757 => x"b9600800", 12758 => x"b8801000",
    12759 => x"f8000027", 12760 => x"b8206000", 12761 => x"b9600800",
    12762 => x"f8001046", 12763 => x"b9800800", 12764 => x"2b9d0004",
    12765 => x"2b8b000c", 12766 => x"2b8c0008", 12767 => x"379c000c",
    12768 => x"c3a00000", 12769 => x"379cffe0", 12770 => x"5b9d0004",
    12771 => x"5b83000c", 12772 => x"3783000c", 12773 => x"5b820008",
    12774 => x"5b840010", 12775 => x"5b850014", 12776 => x"5b860018",
    12777 => x"5b87001c", 12778 => x"5b880020", 12779 => x"f8000013",
    12780 => x"2b9d0004", 12781 => x"379c0020", 12782 => x"c3a00000",
    12783 => x"379cffdc", 12784 => x"5b9d0004", 12785 => x"5b82000c",
    12786 => x"3782000c", 12787 => x"5b810008", 12788 => x"5b830010",
    12789 => x"5b840014", 12790 => x"5b850018", 12791 => x"5b86001c",
    12792 => x"5b870020", 12793 => x"5b880024", 12794 => x"fbffffd3",
    12795 => x"2b9d0004", 12796 => x"379c0024", 12797 => x"c3a00000",
    12798 => x"379cff94", 12799 => x"5b8b0044", 12800 => x"5b8c0040",
    12801 => x"5b8d003c", 12802 => x"5b8e0038", 12803 => x"5b8f0034",
    12804 => x"5b900030", 12805 => x"5b91002c", 12806 => x"5b920028",
    12807 => x"5b930024", 12808 => x"5b940020", 12809 => x"5b95001c",
    12810 => x"5b960018", 12811 => x"5b970014", 12812 => x"5b980010",
    12813 => x"5b99000c", 12814 => x"5b9b0008", 12815 => x"5b9d0004",
    12816 => x"78160001", 12817 => x"b820c800", 12818 => x"b840a000",
    12819 => x"b8209800", 12820 => x"34180025", 12821 => x"34090069",
    12822 => x"34080070", 12823 => x"34070058", 12824 => x"34060063",
    12825 => x"34050064", 12826 => x"341b002a", 12827 => x"340a0030",
    12828 => x"34170010", 12829 => x"37950060", 12830 => x"3ad65620",
    12831 => x"e0000093", 12832 => x"34110001", 12833 => x"34100020",
    12834 => x"340e000a", 12835 => x"44380004", 12836 => x"32610000",
    12837 => x"e0000038", 12838 => x"34100030", 12839 => x"36940001",
    12840 => x"42810000", 12841 => x"4429003c", 12842 => x"5429000d",
    12843 => x"44270037", 12844 => x"54270008", 12845 => x"443b0018",
    12846 => x"543b0004", 12847 => x"44200085", 12848 => x"5c380017",
    12849 => x"e000002b", 12850 => x"5c2a0015", 12851 => x"e3fffff3",
    12852 => x"44260019", 12853 => x"5c250012", 12854 => x"e000002f",
    12855 => x"4428002b", 12856 => x"54280006", 12857 => x"3402006e",
    12858 => x"44220077", 12859 => x"3404006f", 12860 => x"5c24000b",
    12861 => x"e0000022", 12862 => x"34020075", 12863 => x"44220026",
    12864 => x"34040078", 12865 => x"44240021", 12866 => x"34020073",
    12867 => x"5c220004", 12868 => x"e000000e", 12869 => x"286e0000",
    12870 => x"34630004", 12871 => x"3422ffcf", 12872 => x"204200ff",
    12873 => x"34040008", 12874 => x"5444ffdd", 12875 => x"3431ffd0",
    12876 => x"e3ffffdb", 12877 => x"28610000", 12878 => x"34630004",
    12879 => x"32610000", 12880 => x"36730001", 12881 => x"e0000060",
    12882 => x"b8600800", 12883 => x"28210000", 12884 => x"34630004",
    12885 => x"e0000004", 12886 => x"32620000", 12887 => x"34210001",
    12888 => x"36730001", 12889 => x"40220000", 12890 => x"5c40fffc",
    12891 => x"e0000056", 12892 => x"32780000", 12893 => x"36730001",
    12894 => x"e0000053", 12895 => x"3401000a", 12896 => x"45c10004",
    12897 => x"e0000004", 12898 => x"340e0010", 12899 => x"e0000002",
    12900 => x"340e0008", 12901 => x"286d0000", 12902 => x"34720004",
    12903 => x"65c3000a", 12904 => x"01a4001f", 12905 => x"340f0000",
    12906 => x"a0831800", 12907 => x"44600003", 12908 => x"c80d6800",
    12909 => x"340f0001", 12910 => x"340c0010", 12911 => x"e0000019",
    12912 => x"b9a00800", 12913 => x"b9c01000", 12914 => x"5b85004c",
    12915 => x"5b860050", 12916 => x"5b870054", 12917 => x"5b880058",
    12918 => x"5b89005c", 12919 => x"5b8a0048", 12920 => x"f80018fa",
    12921 => x"b6c11800", 12922 => x"40630000", 12923 => x"358cffff",
    12924 => x"b6ac5800", 12925 => x"b9a00800", 12926 => x"31630000",
    12927 => x"b9c01000", 12928 => x"f80018e2", 12929 => x"2b8a0048",
    12930 => x"2b89005c", 12931 => x"2b880058", 12932 => x"2b870054",
    12933 => x"2b860050", 12934 => x"2b85004c", 12935 => x"b8206800",
    12936 => x"7d840000", 12937 => x"7da30000", 12938 => x"a0831800",
    12939 => x"5c60ffe5", 12940 => x"5d970004", 12941 => x"34020030",
    12942 => x"3382006f", 12943 => x"340c000f", 12944 => x"66020020",
    12945 => x"a1e21000", 12946 => x"4440000b", 12947 => x"358cffff",
    12948 => x"b6ac1000", 12949 => x"3403002d", 12950 => x"30430000",
    12951 => x"340f0000", 12952 => x"e0000005", 12953 => x"358cffff",
    12954 => x"b6ac1000", 12955 => x"30500000", 12956 => x"e0000003",
    12957 => x"caf10800", 12958 => x"b42f0800", 12959 => x"4981fffa",
    12960 => x"45e00005", 12961 => x"358cffff", 12962 => x"b6ac0800",
    12963 => x"3402002d", 12964 => x"30220000", 12965 => x"caec1800",
    12966 => x"ba600800", 12967 => x"3404000f", 12968 => x"e0000006",
    12969 => x"b6ac1000", 12970 => x"40420000", 12971 => x"358c0001",
    12972 => x"30220000", 12973 => x"34210001", 12974 => x"4c8cfffb",
    12975 => x"b6639800", 12976 => x"ba401800", 12977 => x"36940001",
    12978 => x"42810000", 12979 => x"5c20ff6d", 12980 => x"ca790800",
    12981 => x"32600000", 12982 => x"2b9d0004", 12983 => x"2b8b0044",
    12984 => x"2b8c0040", 12985 => x"2b8d003c", 12986 => x"2b8e0038",
    12987 => x"2b8f0034", 12988 => x"2b900030", 12989 => x"2b91002c",
    12990 => x"2b920028", 12991 => x"2b930024", 12992 => x"2b940020",
    12993 => x"2b95001c", 12994 => x"2b960018", 12995 => x"2b970014",
    12996 => x"2b980010", 12997 => x"2b99000c", 12998 => x"2b9b0008",
    12999 => x"379c006c", 13000 => x"c3a00000", 13001 => x"78020001",
    13002 => x"14210002", 13003 => x"384292ac", 13004 => x"28420000",
    13005 => x"202100ff", 13006 => x"3c210010", 13007 => x"5841002c",
    13008 => x"28410030", 13009 => x"4c20ffff", 13010 => x"28410030",
    13011 => x"2021ffff", 13012 => x"c3a00000", 13013 => x"14210002",
    13014 => x"78030001", 13015 => x"386392ac", 13016 => x"202100ff",
    13017 => x"28630000", 13018 => x"2042ffff", 13019 => x"78048000",
    13020 => x"3c210010", 13021 => x"b8441000", 13022 => x"b8411000",
    13023 => x"5862002c", 13024 => x"28610030", 13025 => x"4c20ffff",
    13026 => x"c3a00000", 13027 => x"40240002", 13028 => x"40230003",
    13029 => x"78020001", 13030 => x"3c840018", 13031 => x"3c630010",
    13032 => x"384292ac", 13033 => x"b8831800", 13034 => x"40240005",
    13035 => x"28420000", 13036 => x"b8641800", 13037 => x"40240004",
    13038 => x"3c840008", 13039 => x"b8641800", 13040 => x"58430028",
    13041 => x"40230001", 13042 => x"40210000", 13043 => x"3c210008",
    13044 => x"b8610800", 13045 => x"58410024", 13046 => x"c3a00000",
    13047 => x"78020001", 13048 => x"384292ac", 13049 => x"28430000",
    13050 => x"28630028", 13051 => x"30230005", 13052 => x"28430000",
    13053 => x"28630028", 13054 => x"00630008", 13055 => x"30230004",
    13056 => x"28430000", 13057 => x"28630028", 13058 => x"00630010",
    13059 => x"30230003", 13060 => x"28430000", 13061 => x"28630028",
    13062 => x"00630018", 13063 => x"30230002", 13064 => x"28430000",
    13065 => x"28630024", 13066 => x"30230001", 13067 => x"28420000",
    13068 => x"28420024", 13069 => x"00420008", 13070 => x"30220000",
    13071 => x"c3a00000", 13072 => x"379cfff4", 13073 => x"5b8b000c",
    13074 => x"5b8c0008", 13075 => x"5b9d0004", 13076 => x"780b0001",
    13077 => x"b8406000", 13078 => x"396b92ac", 13079 => x"5c200004",
    13080 => x"29610000", 13081 => x"58200000", 13082 => x"e0000022",
    13083 => x"29610000", 13084 => x"58200000", 13085 => x"28220034",
    13086 => x"78010001", 13087 => x"38215634", 13088 => x"fbfffecf",
    13089 => x"f80000be", 13090 => x"29610000", 13091 => x"340200e0",
    13092 => x"58220000", 13093 => x"78010001", 13094 => x"382182c0",
    13095 => x"34020800", 13096 => x"582c0000", 13097 => x"34010000",
    13098 => x"fbffffab", 13099 => x"340100c8", 13100 => x"f8000488",
    13101 => x"34010000", 13102 => x"38028000", 13103 => x"fbffffa6",
    13104 => x"34010000", 13105 => x"34020000", 13106 => x"fbffffa3",
    13107 => x"34010010", 13108 => x"34020000", 13109 => x"fbffffa0",
    13110 => x"7d820000", 13111 => x"34010000", 13112 => x"c8021000",
    13113 => x"20421200", 13114 => x"34420140", 13115 => x"fbffff9a",
    13116 => x"34010000", 13117 => x"2b9d0004", 13118 => x"2b8b000c",
    13119 => x"2b8c0008", 13120 => x"379c000c", 13121 => x"c3a00000",
    13122 => x"379cfff0", 13123 => x"5b8b000c", 13124 => x"5b8c0008",
    13125 => x"5b9d0004", 13126 => x"78020001", 13127 => x"384282c0",
    13128 => x"284b0000", 13129 => x"b8206000", 13130 => x"34010004",
    13131 => x"fbffff7e", 13132 => x"7d6b0000", 13133 => x"0f810012",
    13134 => x"34010004", 13135 => x"c80b5800", 13136 => x"fbffff79",
    13137 => x"216b0020", 13138 => x"0f810012", 13139 => x"356b0004",
    13140 => x"45800004", 13141 => x"34010014", 13142 => x"fbffff73",
    13143 => x"0d810000", 13144 => x"2f810012", 13145 => x"a1610800",
    13146 => x"e42b0800", 13147 => x"2b9d0004", 13148 => x"2b8b000c",
    13149 => x"2b8c0008", 13150 => x"379c0010", 13151 => x"c3a00000",
    13152 => x"379cfffc", 13153 => x"5b9d0004", 13154 => x"34010040",
    13155 => x"fbffff66", 13156 => x"00210004", 13157 => x"2021001f",
    13158 => x"08210320", 13159 => x"2b9d0004", 13160 => x"379c0004",
    13161 => x"c3a00000", 13162 => x"379cfff4", 13163 => x"5b8b000c",
    13164 => x"5b8c0008", 13165 => x"5b9d0004", 13166 => x"78030001",
    13167 => x"38638ec8", 13168 => x"b8405800", 13169 => x"28620000",
    13170 => x"58220000", 13171 => x"78010001", 13172 => x"38218ecc",
    13173 => x"282c0000", 13174 => x"34010040", 13175 => x"fbffff52",
    13176 => x"00210004", 13177 => x"2021001f", 13178 => x"08210320",
    13179 => x"b42c0800", 13180 => x"59610000", 13181 => x"34010000",
    13182 => x"2b9d0004", 13183 => x"2b8b000c", 13184 => x"2b8c0008",
    13185 => x"379c000c", 13186 => x"c3a00000", 13187 => x"379cfffc",
    13188 => x"5b9d0004", 13189 => x"34010040", 13190 => x"fbffff43",
    13191 => x"38220001", 13192 => x"34010040", 13193 => x"fbffff4c",
    13194 => x"34010000", 13195 => x"2b9d0004", 13196 => x"379c0004",
    13197 => x"c3a00000", 13198 => x"379cfffc", 13199 => x"5b9d0004",
    13200 => x"34010040", 13201 => x"fbffff38", 13202 => x"3402fffe",
    13203 => x"a0221000", 13204 => x"34010040", 13205 => x"fbffff40",
    13206 => x"34010000", 13207 => x"2b9d0004", 13208 => x"379c0004",
    13209 => x"c3a00000", 13210 => x"379cfff8", 13211 => x"5b8b0008",
    13212 => x"5b9d0004", 13213 => x"780b0001", 13214 => x"396b92ac",
    13215 => x"29610000", 13216 => x"28220004", 13217 => x"38420010",
    13218 => x"58220004", 13219 => x"34010001", 13220 => x"f8000410",
    13221 => x"29610000", 13222 => x"28210004", 13223 => x"20210020",
    13224 => x"7c210000", 13225 => x"2b9d0004", 13226 => x"2b8b0008",
    13227 => x"379c0008", 13228 => x"c3a00000", 13229 => x"379cfff8",
    13230 => x"5b8b0008", 13231 => x"5b9d0004", 13232 => x"b8205800",
    13233 => x"34010044", 13234 => x"fbffff17", 13235 => x"38220020",
    13236 => x"45600003", 13237 => x"3402ffdf", 13238 => x"a0221000",
    13239 => x"34010044", 13240 => x"fbffff1d", 13241 => x"34010000",
    13242 => x"2b9d0004", 13243 => x"2b8b0008", 13244 => x"379c0008",
    13245 => x"c3a00000", 13246 => x"379cfff8", 13247 => x"5b8b0008",
    13248 => x"5b9d0004", 13249 => x"78020001", 13250 => x"38428f28",
    13251 => x"28420000", 13252 => x"780b0001", 13253 => x"396b92ac",
    13254 => x"59620000", 13255 => x"fbffff1c", 13256 => x"34010001",
    13257 => x"fbffffe4", 13258 => x"78020001", 13259 => x"38425a6c",
    13260 => x"28410000", 13261 => x"78040001", 13262 => x"38845a70",
    13263 => x"58200000", 13264 => x"29610000", 13265 => x"28830000",
    13266 => x"34020003", 13267 => x"58200000", 13268 => x"5822000c",
    13269 => x"58230008", 13270 => x"78030001", 13271 => x"38635a74",
    13272 => x"58220004", 13273 => x"28620000", 13274 => x"5822003c",
    13275 => x"2b9d0004", 13276 => x"2b8b0008", 13277 => x"379c0008",
    13278 => x"c3a00000", 13279 => x"379cffec", 13280 => x"5b8b000c",
    13281 => x"5b8c0008", 13282 => x"5b9d0004", 13283 => x"78010001",
    13284 => x"3821757c", 13285 => x"28220000", 13286 => x"78010001",
    13287 => x"38216fdc", 13288 => x"44400003", 13289 => x"78010001",
    13290 => x"38216fe4", 13291 => x"282b0000", 13292 => x"5d600004",
    13293 => x"78010001", 13294 => x"3821563c", 13295 => x"e0000036",
    13296 => x"78030001", 13297 => x"38635a78", 13298 => x"282c0004",
    13299 => x"29620000", 13300 => x"28610000", 13301 => x"44410011",
    13302 => x"b9600800", 13303 => x"780400ff", 13304 => x"e000000d",
    13305 => x"28230000", 13306 => x"3c660018", 13307 => x"00650018",
    13308 => x"b8c52800", 13309 => x"a0643000", 13310 => x"00c60008",
    13311 => x"2063ff00", 13312 => x"3c630008", 13313 => x"b8a62800",
    13314 => x"b8a31800", 13315 => x"58230000", 13316 => x"34210004",
    13317 => x"5581fff4", 13318 => x"78040001", 13319 => x"38845a78",
    13320 => x"29630000", 13321 => x"28810000", 13322 => x"44610005",
    13323 => x"78010001", 13324 => x"38215654", 13325 => x"fbfffde2",
    13326 => x"e000008c", 13327 => x"78010001", 13328 => x"382182c4",
    13329 => x"28220000", 13330 => x"356b0004", 13331 => x"5c400016",
    13332 => x"29630008", 13333 => x"34021234", 13334 => x"0063000d",
    13335 => x"2063ffff", 13336 => x"5c62000b", 13337 => x"29630010",
    13338 => x"34025678", 13339 => x"0063000d", 13340 => x"2063ffff",
    13341 => x"5c620006", 13342 => x"29630018", 13343 => x"34424444",
    13344 => x"0063000d", 13345 => x"2063ffff", 13346 => x"44620005",
    13347 => x"78010001", 13348 => x"3821567c", 13349 => x"fbfffdca",
    13350 => x"e0000074", 13351 => x"34020001", 13352 => x"58220000",
    13353 => x"37810010", 13354 => x"fbfffecd", 13355 => x"78050001",
    13356 => x"38a55a7c", 13357 => x"28a20000", 13358 => x"29640008",
    13359 => x"29630010", 13360 => x"29610018", 13361 => x"a0822000",
    13362 => x"a0621800", 13363 => x"a0220800", 13364 => x"59640008",
    13365 => x"59630010", 13366 => x"59610018", 13367 => x"43850010",
    13368 => x"43860011", 13369 => x"3ca50008", 13370 => x"b8a62800",
    13371 => x"3ca5000d", 13372 => x"3806cafe", 13373 => x"b8852000",
    13374 => x"59640008", 13375 => x"43840012", 13376 => x"43850013",
    13377 => x"3c840008", 13378 => x"b8852000", 13379 => x"3c84000d",
    13380 => x"34050001", 13381 => x"b8641800", 13382 => x"59630010",
    13383 => x"43830014", 13384 => x"43840015", 13385 => x"3c630008",
    13386 => x"b8641800", 13387 => x"3c63000d", 13388 => x"b8230800",
    13389 => x"78030001", 13390 => x"38635a80", 13391 => x"59610018",
    13392 => x"28640000", 13393 => x"b9600800", 13394 => x"e000000b",
    13395 => x"28230000", 13396 => x"0067000d", 13397 => x"20e7ffff",
    13398 => x"5ce60006", 13399 => x"20670007", 13400 => x"5ce50004",
    13401 => x"a0621800", 13402 => x"b8641800", 13403 => x"58230000",
    13404 => x"34210008", 13405 => x"5581fff6", 13406 => x"78040001",
    13407 => x"38845a7c", 13408 => x"78030001", 13409 => x"b9600800",
    13410 => x"34020000", 13411 => x"34070aaa", 13412 => x"34060007",
    13413 => x"28850000", 13414 => x"3863757c", 13415 => x"e0000010",
    13416 => x"28240000", 13417 => x"0088000d", 13418 => x"2108ffff",
    13419 => x"5d07000b", 13420 => x"00880007", 13421 => x"2108001f",
    13422 => x"5d060008", 13423 => x"a0852000", 13424 => x"58240000",
    13425 => x"28620000", 13426 => x"3c42000d", 13427 => x"b8442000",
    13428 => x"58240000", 13429 => x"b8201000", 13430 => x"34210008",
    13431 => x"5581fff1", 13432 => x"78010001", 13433 => x"382192ac",
    13434 => x"28210000", 13435 => x"34030000", 13436 => x"58200014",
    13437 => x"e000000f", 13438 => x"29640000", 13439 => x"29660004",
    13440 => x"356b0008", 13441 => x"20850fff", 13442 => x"3cc60014",
    13443 => x"0084000c", 13444 => x"58250018", 13445 => x"b8c42000",
    13446 => x"3c840008", 13447 => x"2066003f", 13448 => x"38840040",
    13449 => x"b8862000", 13450 => x"58240014", 13451 => x"34630001",
    13452 => x"558bfff2", 13453 => x"4440000b", 13454 => x"78050001",
    13455 => x"38a55a7c", 13456 => x"28440000", 13457 => x"28a30000",
    13458 => x"78050001", 13459 => x"38a55a84", 13460 => x"a0831800",
    13461 => x"28a40000", 13462 => x"b8641800", 13463 => x"58430000",
    13464 => x"34020080", 13465 => x"58220014", 13466 => x"2b9d0004",
    13467 => x"2b8b000c", 13468 => x"2b8c0008", 13469 => x"379c0014",
    13470 => x"c3a00000", 13471 => x"78030001", 13472 => x"386392a8",
    13473 => x"44400004", 13474 => x"28620000", 13475 => x"58410004",
    13476 => x"c3a00000", 13477 => x"28620000", 13478 => x"58410008",
    13479 => x"c3a00000", 13480 => x"78030001", 13481 => x"386392a8",
    13482 => x"44400004", 13483 => x"28620000", 13484 => x"58410004",
    13485 => x"c3a00000", 13486 => x"28620000", 13487 => x"58410008",
    13488 => x"c3a00000", 13489 => x"3401012c", 13490 => x"34000000",
    13491 => x"3421ffff", 13492 => x"5c20fffe", 13493 => x"c3a00000",
    13494 => x"379cfff8", 13495 => x"5b8b0008", 13496 => x"5b9d0004",
    13497 => x"202100ff", 13498 => x"3c2b0003", 13499 => x"78020001",
    13500 => x"38426fec", 13501 => x"b44b5800", 13502 => x"29610004",
    13503 => x"34020000", 13504 => x"fbffffdf", 13505 => x"fbfffff0",
    13506 => x"29610000", 13507 => x"34020000", 13508 => x"fbffffdb",
    13509 => x"fbffffec", 13510 => x"2b9d0004", 13511 => x"2b8b0008",
    13512 => x"379c0008", 13513 => x"c3a00000", 13514 => x"379cfff8",
    13515 => x"5b8b0008", 13516 => x"5b9d0004", 13517 => x"202100ff",
    13518 => x"3c2b0003", 13519 => x"78020001", 13520 => x"38426fec",
    13521 => x"b44b5800", 13522 => x"29610004", 13523 => x"34020001",
    13524 => x"fbffffcb", 13525 => x"fbffffdc", 13526 => x"29610000",
    13527 => x"34020001", 13528 => x"fbffffc7", 13529 => x"fbffffd8",
    13530 => x"29610004", 13531 => x"34020000", 13532 => x"fbffffc3",
    13533 => x"fbffffd4", 13534 => x"29610000", 13535 => x"34020000",
    13536 => x"fbffffbf", 13537 => x"fbffffd0", 13538 => x"2b9d0004",
    13539 => x"2b8b0008", 13540 => x"379c0008", 13541 => x"c3a00000",
    13542 => x"379cfff8", 13543 => x"5b8b0008", 13544 => x"5b9d0004",
    13545 => x"202100ff", 13546 => x"3c2b0003", 13547 => x"78020001",
    13548 => x"38426fec", 13549 => x"b44b5800", 13550 => x"29610004",
    13551 => x"34020000", 13552 => x"fbffffaf", 13553 => x"fbffffc0",
    13554 => x"29610000", 13555 => x"34020001", 13556 => x"fbffffab",
    13557 => x"fbffffbc", 13558 => x"29610004", 13559 => x"34020001",
    13560 => x"fbffffa7", 13561 => x"fbffffb8", 13562 => x"2b9d0004",
    13563 => x"2b8b0008", 13564 => x"379c0008", 13565 => x"c3a00000",
    13566 => x"379cffec", 13567 => x"5b8b0014", 13568 => x"5b8c0010",
    13569 => x"5b8d000c", 13570 => x"5b8e0008", 13571 => x"5b9d0004",
    13572 => x"202100ff", 13573 => x"78030001", 13574 => x"3c2b0003",
    13575 => x"38636fec", 13576 => x"204e00ff", 13577 => x"340d0008",
    13578 => x"b46b5800", 13579 => x"29610004", 13580 => x"21c20080",
    13581 => x"35adffff", 13582 => x"fbffff91", 13583 => x"fbffffa2",
    13584 => x"29610000", 13585 => x"34020001", 13586 => x"3dce0001",
    13587 => x"fbffff8c", 13588 => x"fbffff9d", 13589 => x"29610000",
    13590 => x"34020000", 13591 => x"21ad00ff", 13592 => x"fbffff87",
    13593 => x"356c0004", 13594 => x"fbffff97", 13595 => x"21ce00ff",
    13596 => x"5da0ffef", 13597 => x"29810000", 13598 => x"34020001",
    13599 => x"fbffff80", 13600 => x"fbffff91", 13601 => x"29610000",
    13602 => x"34020001", 13603 => x"fbffff7c", 13604 => x"fbffff8d",
    13605 => x"78010001", 13606 => x"382192a8", 13607 => x"28210000",
    13608 => x"298d0000", 13609 => x"34020000", 13610 => x"28210004",
    13611 => x"a02d6800", 13612 => x"29610000", 13613 => x"fbffff72",
    13614 => x"fbffff83", 13615 => x"29810000", 13616 => x"34020000",
    13617 => x"fbffff6e", 13618 => x"fbffff7f", 13619 => x"7da10000",
    13620 => x"2b9d0004", 13621 => x"2b8b0014", 13622 => x"2b8c0010",
    13623 => x"2b8d000c", 13624 => x"2b8e0008", 13625 => x"379c0014",
    13626 => x"c3a00000", 13627 => x"379cffe0", 13628 => x"5b8b0020",
    13629 => x"5b8c001c", 13630 => x"5b8d0018", 13631 => x"5b8e0014",
    13632 => x"5b8f0010", 13633 => x"5b90000c", 13634 => x"5b910008",
    13635 => x"5b9d0004", 13636 => x"202100ff", 13637 => x"3c2b0003",
    13638 => x"78040001", 13639 => x"38846fec", 13640 => x"b48b5800",
    13641 => x"29610004", 13642 => x"b8407800", 13643 => x"34020001",
    13644 => x"207000ff", 13645 => x"fbffff52", 13646 => x"fbffff63",
    13647 => x"29610000", 13648 => x"34020000", 13649 => x"780d0001",
    13650 => x"fbffff4d", 13651 => x"340c0000", 13652 => x"fbffff5d",
    13653 => x"340e0000", 13654 => x"39ad92a8", 13655 => x"34110008",
    13656 => x"29610000", 13657 => x"34020001", 13658 => x"3d8c0001",
    13659 => x"fbffff44", 13660 => x"fbffff55", 13661 => x"29a10000",
    13662 => x"29620004", 13663 => x"218c00ff", 13664 => x"28210004",
    13665 => x"a0220800", 13666 => x"44200002", 13667 => x"398c0001",
    13668 => x"29610000", 13669 => x"34020000", 13670 => x"35ce0001",
    13671 => x"fbffff38", 13672 => x"fbffff49", 13673 => x"5dd1ffef",
    13674 => x"46000004", 13675 => x"29610004", 13676 => x"34020001",
    13677 => x"e0000003", 13678 => x"29610004", 13679 => x"34020000",
    13680 => x"fbffff2f", 13681 => x"fbffff40", 13682 => x"29610000",
    13683 => x"34020001", 13684 => x"fbffff2b", 13685 => x"fbffff3c",
    13686 => x"29610000", 13687 => x"34020000", 13688 => x"fbffff27",
    13689 => x"fbffff38", 13690 => x"31ec0000", 13691 => x"2b9d0004",
    13692 => x"2b8b0020", 13693 => x"2b8c001c", 13694 => x"2b8d0018",
    13695 => x"2b8e0014", 13696 => x"2b8f0010", 13697 => x"2b90000c",
    13698 => x"2b910008", 13699 => x"379c0020", 13700 => x"c3a00000",
    13701 => x"379cfff8", 13702 => x"5b8b0008", 13703 => x"5b9d0004",
    13704 => x"202100ff", 13705 => x"3c2b0003", 13706 => x"78020001",
    13707 => x"38426fec", 13708 => x"b44b5800", 13709 => x"29610000",
    13710 => x"34020001", 13711 => x"fbffff10", 13712 => x"fbffff21",
    13713 => x"29610004", 13714 => x"34020001", 13715 => x"fbffff0c",
    13716 => x"fbffff1d", 13717 => x"2b9d0004", 13718 => x"2b8b0008",
    13719 => x"379c0008", 13720 => x"c3a00000", 13721 => x"379cfff4",
    13722 => x"5b8b000c", 13723 => x"5b8c0008", 13724 => x"5b9d0004",
    13725 => x"202b00ff", 13726 => x"b9600800", 13727 => x"204c00ff",
    13728 => x"fbffff16", 13729 => x"3d820001", 13730 => x"b9600800",
    13731 => x"204200fe", 13732 => x"fbffff5a", 13733 => x"b8206000",
    13734 => x"b9600800", 13735 => x"fbffff3f", 13736 => x"65810000",
    13737 => x"2b9d0004", 13738 => x"2b8b000c", 13739 => x"2b8c0008",
    13740 => x"379c000c", 13741 => x"c3a00000", 13742 => x"379cffe8",
    13743 => x"5b8b0018", 13744 => x"5b8c0014", 13745 => x"5b8d0010",
    13746 => x"5b8e000c", 13747 => x"5b8f0008", 13748 => x"5b9d0004",
    13749 => x"780b0001", 13750 => x"396b925c", 13751 => x"296d000c",
    13752 => x"296f0004", 13753 => x"b8206000", 13754 => x"3dad0002",
    13755 => x"c84f0800", 13756 => x"b9a01000", 13757 => x"b8607000",
    13758 => x"f80015b4", 13759 => x"b42f1000", 13760 => x"b5af6800",
    13761 => x"b44e0800", 13762 => x"542d0006", 13763 => x"b9800800",
    13764 => x"b9c01800", 13765 => x"f80015fe", 13766 => x"b8206000",
    13767 => x"e0000009", 13768 => x"c9a26800", 13769 => x"b9a01800",
    13770 => x"b9800800", 13771 => x"f80015f8", 13772 => x"29620004",
    13773 => x"b58d0800", 13774 => x"c9cd1800", 13775 => x"f80015f4",
    13776 => x"b9800800", 13777 => x"2b9d0004", 13778 => x"2b8b0018",
    13779 => x"2b8c0014", 13780 => x"2b8d0010", 13781 => x"2b8e000c",
    13782 => x"2b8f0008", 13783 => x"379c0018", 13784 => x"c3a00000",
    13785 => x"379cffe8", 13786 => x"5b8b0018", 13787 => x"5b8c0014",
    13788 => x"5b8d0010", 13789 => x"5b8e000c", 13790 => x"5b8f0008",
    13791 => x"5b9d0004", 13792 => x"780b0001", 13793 => x"396b925c",
    13794 => x"296f000c", 13795 => x"296e0004", 13796 => x"b8406800",
    13797 => x"3def0002", 13798 => x"c82e0800", 13799 => x"b9e01000",
    13800 => x"f800158a", 13801 => x"b42e6000", 13802 => x"b58d0800",
    13803 => x"b5ee7000", 13804 => x"542e0006", 13805 => x"b9800800",
    13806 => x"34020000", 13807 => x"b9a01800", 13808 => x"f8001651",
    13809 => x"e000000b", 13810 => x"c9cc7000", 13811 => x"34020000",
    13812 => x"b9c01800", 13813 => x"b9800800", 13814 => x"f800164b",
    13815 => x"29610004", 13816 => x"34020000", 13817 => x"c9ae1800",
    13818 => x"f8001647", 13819 => x"b9800800", 13820 => x"2b9d0004",
    13821 => x"2b8b0018", 13822 => x"2b8c0014", 13823 => x"2b8d0010",
    13824 => x"2b8e000c", 13825 => x"2b8f0008", 13826 => x"379c0018",
    13827 => x"c3a00000", 13828 => x"379cfff4", 13829 => x"5b8b000c",
    13830 => x"5b8c0008", 13831 => x"5b9d0004", 13832 => x"780c0001",
    13833 => x"398c92bc", 13834 => x"29810000", 13835 => x"780b0001",
    13836 => x"396b925c", 13837 => x"58200000", 13838 => x"34020200",
    13839 => x"78010001", 13840 => x"382186c8", 13841 => x"5962000c",
    13842 => x"34020800", 13843 => x"59610004", 13844 => x"59610000",
    13845 => x"fbffffc4", 13846 => x"29620004", 13847 => x"29810000",
    13848 => x"58220008", 13849 => x"2962000c", 13850 => x"5822000c",
    13851 => x"34020002", 13852 => x"5822004c", 13853 => x"34020400",
    13854 => x"58220000", 13855 => x"2b9d0004", 13856 => x"2b8b000c",
    13857 => x"2b8c0008", 13858 => x"379c000c", 13859 => x"c3a00000",
    13860 => x"379cfff4", 13861 => x"5b8b000c", 13862 => x"5b8c0008",
    13863 => x"5b9d0004", 13864 => x"780b0001", 13865 => x"396b92bc",
    13866 => x"29630000", 13867 => x"340c0002", 13868 => x"78010001",
    13869 => x"586c0040", 13870 => x"78020001", 13871 => x"586c004c",
    13872 => x"3821925c", 13873 => x"384286c8", 13874 => x"58220004",
    13875 => x"00420002", 13876 => x"34040800", 13877 => x"5824000c",
    13878 => x"344401ff", 13879 => x"3c840010", 13880 => x"2042ffff",
    13881 => x"b8821000", 13882 => x"58620020", 13883 => x"78020001",
    13884 => x"384282c8", 13885 => x"58220014", 13886 => x"34020100",
    13887 => x"5822001c", 13888 => x"58200020", 13889 => x"58200024",
    13890 => x"fbffffc2", 13891 => x"29610000", 13892 => x"582c0044",
    13893 => x"2b9d0004", 13894 => x"2b8b000c", 13895 => x"2b8c0008",
    13896 => x"379c000c", 13897 => x"c3a00000", 13898 => x"379cffc8",
    13899 => x"5b8b0024", 13900 => x"5b8c0020", 13901 => x"5b8d001c",
    13902 => x"5b8e0018", 13903 => x"5b8f0014", 13904 => x"5b900010",
    13905 => x"5b91000c", 13906 => x"5b920008", 13907 => x"5b9d0004",
    13908 => x"b8805800", 13909 => x"78040001", 13910 => x"388492bc",
    13911 => x"b8608000", 13912 => x"28830000", 13913 => x"b8209000",
    13914 => x"b8408800", 13915 => x"2861004c", 13916 => x"340d0000",
    13917 => x"20210002", 13918 => x"4420008b", 13919 => x"780e0001",
    13920 => x"39ce925c", 13921 => x"29c20000", 13922 => x"28440000",
    13923 => x"4804000a", 13924 => x"28610000", 13925 => x"20210200",
    13926 => x"5c200005", 13927 => x"78010001", 13928 => x"382156a4",
    13929 => x"b8801800", 13930 => x"fbfffb85", 13931 => x"fbffff99",
    13932 => x"e000007d", 13933 => x"20810001", 13934 => x"208c0ffe",
    13935 => x"c9816000", 13936 => x"358f0003", 13937 => x"01ef0002",
    13938 => x"78034000", 13939 => x"a0831800", 13940 => x"35ef0001",
    13941 => x"340dffff", 13942 => x"5c600054", 13943 => x"7d610000",
    13944 => x"0084001d", 13945 => x"a0812000", 13946 => x"4483003e",
    13947 => x"b44c1000", 13948 => x"34030004", 13949 => x"37810034",
    13950 => x"fbffff30", 13951 => x"29c30000", 13952 => x"358dfffa",
    13953 => x"358cfffe", 13954 => x"b46c1000", 13955 => x"3781003a",
    13956 => x"34030002", 13957 => x"fbffff29", 13958 => x"78010001",
    13959 => x"38215a88", 13960 => x"282c0000", 13961 => x"37820030",
    13962 => x"37810028", 13963 => x"2b8e0034", 13964 => x"f80004bf",
    13965 => x"78020001", 13966 => x"38425a8c", 13967 => x"28410000",
    13968 => x"a1cc6000", 13969 => x"01ce001c", 13970 => x"502c000e",
    13971 => x"78030001", 13972 => x"38635a90", 13973 => x"2b820030",
    13974 => x"28610000", 13975 => x"54410009", 13976 => x"2b82002c",
    13977 => x"2b810028", 13978 => x"3444ffff", 13979 => x"f4441000",
    13980 => x"3421ffff", 13981 => x"b4410800", 13982 => x"5b810028",
    13983 => x"5b84002c", 13984 => x"78020001", 13985 => x"38425a68",
    13986 => x"28410000", 13987 => x"2b82002c", 13988 => x"2183000f",
    13989 => x"c86e1800", 13990 => x"a0410800", 13991 => x"5961000c",
    13992 => x"6461fff1", 13993 => x"64630001", 13994 => x"59600008",
    13995 => x"b8231800", 13996 => x"44600004", 13997 => x"34010001",
    13998 => x"59610004", 13999 => x"e0000002", 14000 => x"59600004",
    14001 => x"2f81003a", 14002 => x"3d8c0003", 14003 => x"20210800",
    14004 => x"64210000", 14005 => x"596c0010", 14006 => x"31610000",
    14007 => x"b9a06000", 14008 => x"358dfff2", 14009 => x"520d0002",
    14010 => x"ba006800", 14011 => x"780b0001", 14012 => x"396b925c",
    14013 => x"29610024", 14014 => x"29620000", 14015 => x"3403000e",
    14016 => x"34210001", 14017 => x"59610024", 14018 => x"34420004",
    14019 => x"ba400800", 14020 => x"fbfffeea", 14021 => x"29630000",
    14022 => x"ba200800", 14023 => x"34620012", 14024 => x"b9a01800",
    14025 => x"fbfffee5", 14026 => x"780b0001", 14027 => x"396b925c",
    14028 => x"3dee0002", 14029 => x"29610000", 14030 => x"b9c01000",
    14031 => x"fbffff0a", 14032 => x"78030001", 14033 => x"386392bc",
    14034 => x"286c0000", 14035 => x"29610000", 14036 => x"598f0010",
    14037 => x"2962000c", 14038 => x"296f0004", 14039 => x"3c420002",
    14040 => x"c82f0800", 14041 => x"b42e0800", 14042 => x"f8001498",
    14043 => x"b42f0800", 14044 => x"59610000", 14045 => x"29820010",
    14046 => x"28210000", 14047 => x"4801000a", 14048 => x"29810000",
    14049 => x"20210200", 14050 => x"44200002", 14051 => x"fbffff21",
    14052 => x"78010001", 14053 => x"382192bc", 14054 => x"28210000",
    14055 => x"34020002", 14056 => x"5822004c", 14057 => x"b9a00800",
    14058 => x"2b9d0004", 14059 => x"2b8b0024", 14060 => x"2b8c0020",
    14061 => x"2b8d001c", 14062 => x"2b8e0018", 14063 => x"2b8f0014",
    14064 => x"2b900010", 14065 => x"2b91000c", 14066 => x"2b920008",
    14067 => x"379c0038", 14068 => x"c3a00000", 14069 => x"379cffd4",
    14070 => x"5b8b0020", 14071 => x"5b8c001c", 14072 => x"5b8d0018",
    14073 => x"5b8e0014", 14074 => x"5b8f0010", 14075 => x"5b90000c",
    14076 => x"5b910008", 14077 => x"5b9d0004", 14078 => x"780b0001",
    14079 => x"78050001", 14080 => x"396b925c", 14081 => x"38a592bc",
    14082 => x"b8208000", 14083 => x"34010100", 14084 => x"5961001c",
    14085 => x"59610018", 14086 => x"b8806000", 14087 => x"28a10000",
    14088 => x"78040001", 14089 => x"388482c8", 14090 => x"2e0e000c",
    14091 => x"59640014", 14092 => x"59640010", 14093 => x"58240004",
    14094 => x"38018100", 14095 => x"fdc17000", 14096 => x"3401fffc",
    14097 => x"c80e7000", 14098 => x"a1c17000", 14099 => x"35ce0012",
    14100 => x"b5c36800", 14101 => x"b8800800", 14102 => x"b8408800",
    14103 => x"b8607800", 14104 => x"34020000", 14105 => x"35a30004",
    14106 => x"f8001527", 14107 => x"29610010", 14108 => x"b9c01800",
    14109 => x"ba001000", 14110 => x"34210004", 14111 => x"f80014a4",
    14112 => x"29610010", 14113 => x"35ce0004", 14114 => x"ba201000",
    14115 => x"b42e0800", 14116 => x"b9e01800", 14117 => x"f800149e",
    14118 => x"3401003b", 14119 => x"502d0002", 14120 => x"e0000002",
    14121 => x"340d003c", 14122 => x"35a30001", 14123 => x"7d810000",
    14124 => x"00630001", 14125 => x"3c21001e", 14126 => x"78048000",
    14127 => x"b8642000", 14128 => x"b8812000", 14129 => x"78010001",
    14130 => x"3821925c", 14131 => x"28220010", 14132 => x"3c630002",
    14133 => x"78010001", 14134 => x"58440000", 14135 => x"382192bc",
    14136 => x"b4431000", 14137 => x"58400000", 14138 => x"28220000",
    14139 => x"340b0000", 14140 => x"b8207800", 14141 => x"28430000",
    14142 => x"341003e8", 14143 => x"38630001", 14144 => x"58430000",
    14145 => x"29e10000", 14146 => x"282e0000", 14147 => x"21c10002",
    14148 => x"5c200009", 14149 => x"34010001", 14150 => x"356b0001",
    14151 => x"f800006d", 14152 => x"5d70fff9", 14153 => x"78010001",
    14154 => x"382156c4", 14155 => x"b9c01000", 14156 => x"fbfffaa3",
    14157 => x"4580003e", 14158 => x"780b0001", 14159 => x"340e0000",
    14160 => x"396b92bc", 14161 => x"340f0064", 14162 => x"29610000",
    14163 => x"28220000", 14164 => x"20420800", 14165 => x"5c40000a",
    14166 => x"34010001", 14167 => x"35ce0001", 14168 => x"f800005c",
    14169 => x"5dcffff9", 14170 => x"78010001", 14171 => x"382156f4",
    14172 => x"fbfffa93", 14173 => x"340e0000", 14174 => x"e0000003",
    14175 => x"282e0014", 14176 => x"21ce0001", 14177 => x"78010001",
    14178 => x"382192bc", 14179 => x"28210000", 14180 => x"78020001",
    14181 => x"38425a88", 14182 => x"282b0018", 14183 => x"28210014",
    14184 => x"28410000", 14185 => x"3782002c", 14186 => x"a1615800",
    14187 => x"37810024", 14188 => x"f80003df", 14189 => x"78030001",
    14190 => x"38635a8c", 14191 => x"28610000", 14192 => x"502b000e",
    14193 => x"78030001", 14194 => x"38635a90", 14195 => x"2b82002c",
    14196 => x"28610000", 14197 => x"54410009", 14198 => x"2b830028",
    14199 => x"2b820024", 14200 => x"3461ffff", 14201 => x"f4611800",
    14202 => x"3442ffff", 14203 => x"b4621000", 14204 => x"5b820024",
    14205 => x"5b810028", 14206 => x"2b810024", 14207 => x"318e0000",
    14208 => x"3d6b0003", 14209 => x"59810008", 14210 => x"2b810028",
    14211 => x"59800004", 14212 => x"598b0010", 14213 => x"5981000c",
    14214 => x"78010001", 14215 => x"3821925c", 14216 => x"28220020",
    14217 => x"34420001", 14218 => x"58220020", 14219 => x"b9a00800",
    14220 => x"2b9d0004", 14221 => x"2b8b0020", 14222 => x"2b8c001c",
    14223 => x"2b8d0018", 14224 => x"2b8e0014", 14225 => x"2b8f0010",
    14226 => x"2b90000c", 14227 => x"2b910008", 14228 => x"379c002c",
    14229 => x"c3a00000", 14230 => x"78030001", 14231 => x"3863925c",
    14232 => x"28640020", 14233 => x"58240000", 14234 => x"28610024",
    14235 => x"58410000", 14236 => x"c3a00000", 14237 => x"78020001",
    14238 => x"384292c0", 14239 => x"28420000", 14240 => x"78030001",
    14241 => x"386392a8", 14242 => x"58620000", 14243 => x"44200005",
    14244 => x"28430010", 14245 => x"78018000", 14246 => x"b8610800",
    14247 => x"e0000006", 14248 => x"78040001", 14249 => x"38845a68",
    14250 => x"28430010", 14251 => x"28810000", 14252 => x"a0610800",
    14253 => x"58410010", 14254 => x"c3a00000", 14255 => x"78010001",
    14256 => x"382192a8", 14257 => x"28210000", 14258 => x"28210014",
    14259 => x"c3a00000", 14260 => x"78020001", 14261 => x"384292a8",
    14262 => x"28420000", 14263 => x"28430014", 14264 => x"b4230800",
    14265 => x"28430014", 14266 => x"c8611800", 14267 => x"4803fffe",
    14268 => x"c3a00000", 14269 => x"78010001", 14270 => x"382192a8",
    14271 => x"28210000", 14272 => x"28210004", 14273 => x"20210080",
    14274 => x"64210000", 14275 => x"c3a00000", 14276 => x"379cffe0",
    14277 => x"5b8b001c", 14278 => x"5b8c0018", 14279 => x"5b8d0014",
    14280 => x"5b8e0010", 14281 => x"5b8f000c", 14282 => x"5b900008",
    14283 => x"5b9d0004", 14284 => x"b8208000", 14285 => x"34010001",
    14286 => x"fbfffdb7", 14287 => x"34010001", 14288 => x"fbfffce6",
    14289 => x"340200a0", 14290 => x"34010001", 14291 => x"fbfffd2b",
    14292 => x"34020000", 14293 => x"34010001", 14294 => x"fbfffd28",
    14295 => x"34010001", 14296 => x"fbfffcf2", 14297 => x"340200a1",
    14298 => x"34010001", 14299 => x"fbfffd23", 14300 => x"378d0023",
    14301 => x"b9a01000", 14302 => x"34030001", 14303 => x"34010001",
    14304 => x"fbfffd5b", 14305 => x"34010001", 14306 => x"fbfffd04",
    14307 => x"34010001", 14308 => x"438c0023", 14309 => x"fbfffcd1",
    14310 => x"34010001", 14311 => x"340200a1", 14312 => x"fbfffd16",
    14313 => x"340bffd9", 14314 => x"340f000f", 14315 => x"340e0017",
    14316 => x"34030000", 14317 => x"34010001", 14318 => x"b9a01000",
    14319 => x"fbfffd4c", 14320 => x"43830023", 14321 => x"b5836000",
    14322 => x"218c00ff", 14323 => x"556f0003", 14324 => x"b60b0800",
    14325 => x"30230000", 14326 => x"356b0001", 14327 => x"5d6efff5",
    14328 => x"37820023", 14329 => x"34030001", 14330 => x"34010001",
    14331 => x"fbfffd40", 14332 => x"34010001", 14333 => x"fbfffce9",
    14334 => x"43810023", 14335 => x"fc2c6000", 14336 => x"c80c0800",
    14337 => x"2b9d0004", 14338 => x"2b8b001c", 14339 => x"2b8c0018",
    14340 => x"2b8d0014", 14341 => x"2b8e0010", 14342 => x"2b8f000c",
    14343 => x"2b900008", 14344 => x"379c0020", 14345 => x"c3a00000",
    14346 => x"379cffd0", 14347 => x"5b8b0010", 14348 => x"5b8c000c",
    14349 => x"5b8d0008", 14350 => x"5b9d0004", 14351 => x"780b0001",
    14352 => x"396b8f34", 14353 => x"31600000", 14354 => x"fbffffab",
    14355 => x"3403ffed", 14356 => x"44200023", 14357 => x"b9600800",
    14358 => x"fbffffae", 14359 => x"b8206000", 14360 => x"3403fffb",
    14361 => x"5c20001e", 14362 => x"378d0014", 14363 => x"b9601000",
    14364 => x"34030010", 14365 => x"b9a00800", 14366 => x"f8001555",
    14367 => x"b9a00800", 14368 => x"f80004c3", 14369 => x"78020001",
    14370 => x"38428ed0", 14371 => x"5c2c0005", 14372 => x"34010001",
    14373 => x"58410000", 14374 => x"3403fffa", 14375 => x"e0000010",
    14376 => x"2b830028", 14377 => x"78010001", 14378 => x"38218ec8",
    14379 => x"58230000", 14380 => x"2b83002c", 14381 => x"78010001",
    14382 => x"38218ecc", 14383 => x"58230000", 14384 => x"2b830024",
    14385 => x"78010001", 14386 => x"38216ffc", 14387 => x"58230000",
    14388 => x"34010002", 14389 => x"58410000", 14390 => x"34030000",
    14391 => x"b8600800", 14392 => x"2b9d0004", 14393 => x"2b8b0010",
    14394 => x"2b8c000c", 14395 => x"2b8d0008", 14396 => x"379c0030",
    14397 => x"c3a00000", 14398 => x"379cffe0", 14399 => x"5b9b0008",
    14400 => x"341b0020", 14401 => x"b77cd800", 14402 => x"5b8b0020",
    14403 => x"5b8c001c", 14404 => x"5b8d0018", 14405 => x"5b8e0014",
    14406 => x"5b8f0010", 14407 => x"5b90000c", 14408 => x"5b9d0004",
    14409 => x"780b0001", 14410 => x"780c0001", 14411 => x"bb807800",
    14412 => x"34020001", 14413 => x"396b70f0", 14414 => x"398c5724",
    14415 => x"e0000012", 14416 => x"bb808000", 14417 => x"379cffe4",
    14418 => x"378e000b", 14419 => x"01ce0003", 14420 => x"35a2002c",
    14421 => x"3dce0003", 14422 => x"34030014", 14423 => x"b9c00800",
    14424 => x"f800136b", 14425 => x"31c00013", 14426 => x"29a20020",
    14427 => x"29630074", 14428 => x"b9800800", 14429 => x"b9c02000",
    14430 => x"fbfff991", 14431 => x"34020000", 14432 => x"ba00e000",
    14433 => x"b9600800", 14434 => x"f80011ca", 14435 => x"b8206800",
    14436 => x"5c20ffec", 14437 => x"b9e0e000", 14438 => x"2b9d0004",
    14439 => x"2b8b0020", 14440 => x"2b8c001c", 14441 => x"2b8d0018",
    14442 => x"2b8e0014", 14443 => x"2b8f0010", 14444 => x"2b90000c",
    14445 => x"2b9b0008", 14446 => x"379c0020", 14447 => x"c3a00000",
    14448 => x"379cffec", 14449 => x"5b8b0014", 14450 => x"5b8c0010",
    14451 => x"5b8d000c", 14452 => x"5b8e0008", 14453 => x"5b9d0004",
    14454 => x"780b0001", 14455 => x"396b8ed4", 14456 => x"29610000",
    14457 => x"5c200007", 14458 => x"78010001", 14459 => x"382170f0",
    14460 => x"f800118e", 14461 => x"29610000", 14462 => x"34210001",
    14463 => x"59610000", 14464 => x"780b0001", 14465 => x"396b7000",
    14466 => x"780c0001", 14467 => x"356d00f0", 14468 => x"398c70f0",
    14469 => x"e0000009", 14470 => x"29620008", 14471 => x"2963000c",
    14472 => x"29640010", 14473 => x"296e0000", 14474 => x"b9800800",
    14475 => x"f8001253", 14476 => x"59c10000", 14477 => x"356b0018",
    14478 => x"5d6dfff8", 14479 => x"2b9d0004", 14480 => x"2b8b0014",
    14481 => x"2b8c0010", 14482 => x"2b8d000c", 14483 => x"2b8e0008",
    14484 => x"379c0014", 14485 => x"c3a00000", 14486 => x"379cfff4",
    14487 => x"5b8b000c", 14488 => x"5b8c0008", 14489 => x"5b9d0004",
    14490 => x"34020000", 14491 => x"b8206000", 14492 => x"f8000482",
    14493 => x"b8205800", 14494 => x"4c200005", 14495 => x"78010001",
    14496 => x"3821574c", 14497 => x"b9601000", 14498 => x"e0000004",
    14499 => x"29820000", 14500 => x"78010001", 14501 => x"38215778",
    14502 => x"fbfff949", 14503 => x"b9600800", 14504 => x"2b9d0004",
    14505 => x"2b8b000c", 14506 => x"2b8c0008", 14507 => x"379c000c",
    14508 => x"c3a00000", 14509 => x"379cfffc", 14510 => x"5b9d0004",
    14511 => x"78010001", 14512 => x"38218ed8", 14513 => x"58200000",
    14514 => x"78020001", 14515 => x"78010001", 14516 => x"38218eec",
    14517 => x"38428edc", 14518 => x"3403ffff", 14519 => x"58230000",
    14520 => x"58430000", 14521 => x"58200008", 14522 => x"58400008",
    14523 => x"58400004", 14524 => x"58200004", 14525 => x"5840000c",
    14526 => x"5820000c", 14527 => x"34020000", 14528 => x"34010000",
    14529 => x"f8000f41", 14530 => x"2b9d0004", 14531 => x"379c0004",
    14532 => x"c3a00000", 14533 => x"379cfff4", 14534 => x"5b8b000c",
    14535 => x"5b8c0008", 14536 => x"5b9d0004", 14537 => x"b8206000",
    14538 => x"34010000", 14539 => x"f8000fe0", 14540 => x"b8205800",
    14541 => x"34020000", 14542 => x"5c200081", 14543 => x"fbfffacb",
    14544 => x"78030001", 14545 => x"38638edc", 14546 => x"28650008",
    14547 => x"78020001", 14548 => x"38428ed8", 14549 => x"b8202000",
    14550 => x"28420000", 14551 => x"44ab0004", 14552 => x"34010001",
    14553 => x"5ca1001d", 14554 => x"e0000010", 14555 => x"34010001",
    14556 => x"44810005", 14557 => x"28610004", 14558 => x"34210001",
    14559 => x"58610004", 14560 => x"e0000002", 14561 => x"58600004",
    14562 => x"78030001", 14563 => x"38638edc", 14564 => x"28650004",
    14565 => x"34010004", 14566 => x"4c250010", 14567 => x"34010001",
    14568 => x"58610008", 14569 => x"e0000002", 14570 => x"44850003",
    14571 => x"58600004", 14572 => x"e000000a", 14573 => x"28650004",
    14574 => x"34010004", 14575 => x"34a50001", 14576 => x"58650004",
    14577 => x"4c250005", 14578 => x"34010002", 14579 => x"58610008",
    14580 => x"3441fe0c", 14581 => x"5861000c", 14582 => x"78030001",
    14583 => x"38638eec", 14584 => x"28650008", 14585 => x"44a00004",
    14586 => x"34010001", 14587 => x"5ca1001c", 14588 => x"e000000f",
    14589 => x"44850005", 14590 => x"28610004", 14591 => x"34210001",
    14592 => x"58610004", 14593 => x"e0000002", 14594 => x"58600004",
    14595 => x"78030001", 14596 => x"38638eec", 14597 => x"28640004",
    14598 => x"34010004", 14599 => x"4c240010", 14600 => x"34010001",
    14601 => x"58610008", 14602 => x"e0000002", 14603 => x"44800003",
    14604 => x"58600004", 14605 => x"e000000a", 14606 => x"28640004",
    14607 => x"34010004", 14608 => x"34840001", 14609 => x"58640004",
    14610 => x"4c240005", 14611 => x"34010002", 14612 => x"58610008",
    14613 => x"3441fe0c", 14614 => x"5861000c", 14615 => x"3401251b",
    14616 => x"4c220030", 14617 => x"78020001", 14618 => x"38428edc",
    14619 => x"28440008", 14620 => x"34010002", 14621 => x"3402ffff",
    14622 => x"5c810031", 14623 => x"78030001", 14624 => x"38638eec",
    14625 => x"28610008", 14626 => x"5c24002d", 14627 => x"2862000c",
    14628 => x"34011f3f", 14629 => x"e0000002", 14630 => x"3442e0c0",
    14631 => x"4841ffff", 14632 => x"78030001", 14633 => x"38638eec",
    14634 => x"5862000c", 14635 => x"78030001", 14636 => x"38638edc",
    14637 => x"2863000c", 14638 => x"34011f3f", 14639 => x"e0000002",
    14640 => x"3463e0c0", 14641 => x"4861ffff", 14642 => x"78040001",
    14643 => x"38848edc", 14644 => x"5883000c", 14645 => x"4c620003",
    14646 => x"3444f060", 14647 => x"e0000004", 14648 => x"34040000",
    14649 => x"4c430002", 14650 => x"34440fa0", 14651 => x"b4831800",
    14652 => x"0062001f", 14653 => x"b4431800", 14654 => x"14620001",
    14655 => x"4c400003", 14656 => x"34421f40", 14657 => x"e0000004",
    14658 => x"34011f3f", 14659 => x"4c220002", 14660 => x"3442e0c0",
    14661 => x"59820000", 14662 => x"34020001", 14663 => x"e0000008",
    14664 => x"78010001", 14665 => x"34420064", 14666 => x"38218ed8",
    14667 => x"58220000", 14668 => x"34010000", 14669 => x"f8000eb5",
    14670 => x"34020000", 14671 => x"b8400800", 14672 => x"2b9d0004",
    14673 => x"2b8b000c", 14674 => x"2b8c0008", 14675 => x"379c000c",
    14676 => x"c3a00000", 14677 => x"379cfff8", 14678 => x"5b8b0008",
    14679 => x"5b9d0004", 14680 => x"78020001", 14681 => x"b8205800",
    14682 => x"b8400800", 14683 => x"38215798", 14684 => x"fbfff893",
    14685 => x"e0000003", 14686 => x"34010064", 14687 => x"fbfffe55",
    14688 => x"34010000", 14689 => x"fbfff9e1", 14690 => x"4420fffc",
    14691 => x"34010003", 14692 => x"34020000", 14693 => x"34030001",
    14694 => x"f8000dc1", 14695 => x"78020001", 14696 => x"b8400800",
    14697 => x"382157b0", 14698 => x"fbfff885", 14699 => x"e0000003",
    14700 => x"34010064", 14701 => x"fbfffe47", 14702 => x"34010000",
    14703 => x"f8000e82", 14704 => x"4420fffc", 14705 => x"78020001",
    14706 => x"b8400800", 14707 => x"38214d20", 14708 => x"fbfff87b",
    14709 => x"78020001", 14710 => x"b8400800", 14711 => x"382157c0",
    14712 => x"fbfff877", 14713 => x"fbffff34", 14714 => x"b9600800",
    14715 => x"fbffff4a", 14716 => x"4420fffe", 14717 => x"2b9d0004",
    14718 => x"2b8b0008", 14719 => x"379c0008", 14720 => x"c3a00000",
    14721 => x"379cfff0", 14722 => x"5b8b000c", 14723 => x"5b8c0008",
    14724 => x"5b9d0004", 14725 => x"b8405800", 14726 => x"34020003",
    14727 => x"5c220020", 14728 => x"fbffff25", 14729 => x"b9600800",
    14730 => x"fbffff3b", 14731 => x"4420fffe", 14732 => x"4c200002",
    14733 => x"e000001a", 14734 => x"37810010", 14735 => x"34020000",
    14736 => x"f800038e", 14737 => x"b8206000", 14738 => x"48010007",
    14739 => x"29620000", 14740 => x"2b810010", 14741 => x"3443ff38",
    14742 => x"54610003", 14743 => x"344200c8", 14744 => x"50410012",
    14745 => x"34020001", 14746 => x"b9600800", 14747 => x"f8000383",
    14748 => x"78030001", 14749 => x"b8206000", 14750 => x"29620000",
    14751 => x"386357e8", 14752 => x"4c200003", 14753 => x"78030001",
    14754 => x"386357e0", 14755 => x"78010001", 14756 => x"382157f0",
    14757 => x"fbfff84a", 14758 => x"e0000004", 14759 => x"b9600800",
    14760 => x"fbfffeee", 14761 => x"b8206000", 14762 => x"29610000",
    14763 => x"fbffef83", 14764 => x"b9800800", 14765 => x"2b9d0004",
    14766 => x"2b8b000c", 14767 => x"2b8c0008", 14768 => x"379c0010",
    14769 => x"c3a00000", 14770 => x"379cfffc", 14771 => x"5b9d0004",
    14772 => x"34010800", 14773 => x"34020001", 14774 => x"fbfffaf2",
    14775 => x"34010400", 14776 => x"34020000", 14777 => x"fbfffaef",
    14778 => x"34011000", 14779 => x"34020000", 14780 => x"fbfffaec",
    14781 => x"2b9d0004", 14782 => x"379c0004", 14783 => x"c3a00000",
    14784 => x"78010001", 14785 => x"3821929c", 14786 => x"28220000",
    14787 => x"78010001", 14788 => x"38219284", 14789 => x"58220000",
    14790 => x"34010001", 14791 => x"58410000", 14792 => x"c3a00000",
    14793 => x"78010001", 14794 => x"38219284", 14795 => x"28210000",
    14796 => x"34020102", 14797 => x"58220000", 14798 => x"c3a00000",
    14799 => x"379cfff8", 14800 => x"5b8b0008", 14801 => x"5b9d0004",
    14802 => x"780b0001", 14803 => x"396b9284", 14804 => x"29610000",
    14805 => x"28220004", 14806 => x"78010001", 14807 => x"38214e9c",
    14808 => x"fbfff817", 14809 => x"29610000", 14810 => x"34020400",
    14811 => x"58220000", 14812 => x"2b9d0004", 14813 => x"2b8b0008",
    14814 => x"379c0008", 14815 => x"c3a00000", 14816 => x"40230000",
    14817 => x"78020001", 14818 => x"40240001", 14819 => x"384292b0",
    14820 => x"28420000", 14821 => x"3c630008", 14822 => x"b8831800",
    14823 => x"58430010", 14824 => x"40240002", 14825 => x"40230003",
    14826 => x"3c840018", 14827 => x"3c630010", 14828 => x"b8832000",
    14829 => x"40230005", 14830 => x"b8832000", 14831 => x"40230004",
    14832 => x"3c630008", 14833 => x"b8830800", 14834 => x"58410014",
    14835 => x"c3a00000", 14836 => x"40240000", 14837 => x"40230003",
    14838 => x"78020001", 14839 => x"3c840018", 14840 => x"384292b0",
    14841 => x"b8642000", 14842 => x"40230001", 14843 => x"28420000",
    14844 => x"3c630010", 14845 => x"b8832000", 14846 => x"40230002",
    14847 => x"3c630008", 14848 => x"b8832000", 14849 => x"3403ff00",
    14850 => x"58440018", 14851 => x"a0832000", 14852 => x"34840001",
    14853 => x"5844001c", 14854 => x"58430020", 14855 => x"3804ea61",
    14856 => x"3803ea60", 14857 => x"58430024", 14858 => x"58440028",
    14859 => x"40210003", 14860 => x"b4231800", 14861 => x"5843002c",
    14862 => x"78030001", 14863 => x"38635a94", 14864 => x"28610000",
    14865 => x"78030001", 14866 => x"38635a98", 14867 => x"58410030",
    14868 => x"38018cae", 14869 => x"58410034", 14870 => x"28610000",
    14871 => x"58410038", 14872 => x"34011f40", 14873 => x"5841003c",
    14874 => x"c3a00000", 14875 => x"379cfff4", 14876 => x"5b8b000c",
    14877 => x"5b8c0008", 14878 => x"5b9d0004", 14879 => x"780b0001",
    14880 => x"780c0001", 14881 => x"396b7418", 14882 => x"398c7424",
    14883 => x"e0000005", 14884 => x"29620000", 14885 => x"b9600800",
    14886 => x"356b000c", 14887 => x"d8400000", 14888 => x"558bfffc",
    14889 => x"2b9d0004", 14890 => x"2b8b000c", 14891 => x"2b8c0008",
    14892 => x"379c000c", 14893 => x"c3a00000", 14894 => x"379cfff0",
    14895 => x"5b8b0010", 14896 => x"5b8c000c", 14897 => x"5b8d0008",
    14898 => x"5b9d0004", 14899 => x"780b0001", 14900 => x"780d0001",
    14901 => x"340c0000", 14902 => x"396b7418", 14903 => x"39ad7424",
    14904 => x"e0000006", 14905 => x"29620000", 14906 => x"b9600800",
    14907 => x"356b000c", 14908 => x"d8400000", 14909 => x"b5816000",
    14910 => x"55abfffb", 14911 => x"69810000", 14912 => x"2b9d0004",
    14913 => x"2b8b0010", 14914 => x"2b8c000c", 14915 => x"2b8d0008",
    14916 => x"379c0010", 14917 => x"c3a00000", 14918 => x"379cffec",
    14919 => x"5b8b0014", 14920 => x"5b8c0010", 14921 => x"5b8d000c",
    14922 => x"5b8e0008", 14923 => x"5b9d0004", 14924 => x"780b0001",
    14925 => x"780d0001", 14926 => x"b8207000", 14927 => x"396b7418",
    14928 => x"39ad7424", 14929 => x"e000000c", 14930 => x"296c0008",
    14931 => x"e0000007", 14932 => x"b9c01000", 14933 => x"f800124e",
    14934 => x"5c200003", 14935 => x"29810004", 14936 => x"e0000007",
    14937 => x"358c0008", 14938 => x"29810000", 14939 => x"5c20fff9",
    14940 => x"356b000c", 14941 => x"55abfff5", 14942 => x"78018000",
    14943 => x"2b9d0004", 14944 => x"2b8b0014", 14945 => x"2b8c0010",
    14946 => x"2b8d000c", 14947 => x"2b8e0008", 14948 => x"379c0014",
    14949 => x"c3a00000", 14950 => x"b8201800", 14951 => x"5c200008",
    14952 => x"78010001", 14953 => x"78020001", 14954 => x"38217418",
    14955 => x"38427424", 14956 => x"44220003", 14957 => x"28210008",
    14958 => x"c3a00000", 14959 => x"28620008", 14960 => x"34610008",
    14961 => x"5c400016", 14962 => x"78020001", 14963 => x"78040001",
    14964 => x"38427418", 14965 => x"38847424", 14966 => x"e000000f",
    14967 => x"28410008", 14968 => x"e000000a", 14969 => x"5c230008",
    14970 => x"78030001", 14971 => x"3442000c", 14972 => x"38637424",
    14973 => x"34010000", 14974 => x"50430009", 14975 => x"28410008",
    14976 => x"c3a00000", 14977 => x"34210008", 14978 => x"28250000",
    14979 => x"5ca0fff6", 14980 => x"3442000c", 14981 => x"5482fff2",
    14982 => x"34010000", 14983 => x"c3a00000", 14984 => x"379cffc8",
    14985 => x"5b8b0038", 14986 => x"5b8c0034", 14987 => x"5b8d0030",
    14988 => x"5b8e002c", 14989 => x"5b8f0028", 14990 => x"5b900024",
    14991 => x"5b910020", 14992 => x"5b92001c", 14993 => x"5b930018",
    14994 => x"5b940014", 14995 => x"5b950010", 14996 => x"5b96000c",
    14997 => x"5b970008", 14998 => x"5b9d0004", 14999 => x"b8207000",
    15000 => x"34010000", 15001 => x"b840b800", 15002 => x"78140001",
    15003 => x"fbffffcb", 15004 => x"78130001", 15005 => x"78120001",
    15006 => x"78110001", 15007 => x"78100001", 15008 => x"780f0001",
    15009 => x"b8206800", 15010 => x"34150000", 15011 => x"340b0000",
    15012 => x"3a945a24", 15013 => x"3a734e44", 15014 => x"3a52581c",
    15015 => x"78168000", 15016 => x"3a3155f8", 15017 => x"3a10469c",
    15018 => x"39ef55f0", 15019 => x"e0000028", 15020 => x"3562000f",
    15021 => x"b5cb0800", 15022 => x"4ae20006", 15023 => x"78020001",
    15024 => x"38425814", 15025 => x"fbfff730", 15026 => x"b5615800",
    15027 => x"e0000021", 15028 => x"29ac0004", 15029 => x"ba801800",
    15030 => x"46a00002", 15031 => x"ba601800", 15032 => x"29a40000",
    15033 => x"ba401000", 15034 => x"fbfff727", 15035 => x"b42b5800",
    15036 => x"5d960005", 15037 => x"b5cb0800", 15038 => x"b9e01000",
    15039 => x"fbfff722", 15040 => x"e000000e", 15041 => x"4d800006",
    15042 => x"b5cb0800", 15043 => x"ba001000", 15044 => x"fbfff71d",
    15045 => x"c80c6000", 15046 => x"b5615800", 15047 => x"2184ffff",
    15048 => x"08842710", 15049 => x"15830010", 15050 => x"b5cb0800",
    15051 => x"00840010", 15052 => x"ba201000", 15053 => x"fbfff714",
    15054 => x"b42b5800", 15055 => x"b9a00800", 15056 => x"fbffff96",
    15057 => x"b8206800", 15058 => x"36b50001", 15059 => x"5da0ffd9",
    15060 => x"b9600800", 15061 => x"2b9d0004", 15062 => x"2b8b0038",
    15063 => x"2b8c0034", 15064 => x"2b8d0030", 15065 => x"2b8e002c",
    15066 => x"2b8f0028", 15067 => x"2b900024", 15068 => x"2b910020",
    15069 => x"2b92001c", 15070 => x"2b930018", 15071 => x"2b940014",
    15072 => x"2b950010", 15073 => x"2b96000c", 15074 => x"2b970008",
    15075 => x"379c0038", 15076 => x"c3a00000", 15077 => x"379cffa8",
    15078 => x"5b8b0008", 15079 => x"5b9d0004", 15080 => x"378b000c",
    15081 => x"b9600800", 15082 => x"34020050", 15083 => x"fbffff9d",
    15084 => x"78010001", 15085 => x"b9601000", 15086 => x"38214860",
    15087 => x"fbfff700", 15088 => x"34010000", 15089 => x"2b9d0004",
    15090 => x"2b8b0008", 15091 => x"379c0058", 15092 => x"c3a00000",
    15093 => x"78010001", 15094 => x"38218f48", 15095 => x"28210000",
    15096 => x"28220008", 15097 => x"2821000c", 15098 => x"202100ff",
    15099 => x"c3a00000", 15100 => x"78010001", 15101 => x"78030001",
    15102 => x"38635a9c", 15103 => x"38218f48", 15104 => x"28210000",
    15105 => x"28620000", 15106 => x"78040001", 15107 => x"38845aa0",
    15108 => x"58220000", 15109 => x"58200014", 15110 => x"28830000",
    15111 => x"58200018", 15112 => x"58200010", 15113 => x"58230000",
    15114 => x"58220000", 15115 => x"5820001c", 15116 => x"c3a00000",
    15117 => x"78040001", 15118 => x"34050002", 15119 => x"38848f48",
    15120 => x"5c25000e", 15121 => x"28810000", 15122 => x"1444001f",
    15123 => x"20840007", 15124 => x"b4831800", 15125 => x"f4832000",
    15126 => x"00630003", 15127 => x"b4821000", 15128 => x"3c42001d",
    15129 => x"58200014", 15130 => x"58200018", 15131 => x"b8431800",
    15132 => x"58230010", 15133 => x"e0000006", 15134 => x"28810000",
    15135 => x"204200ff", 15136 => x"58230014", 15137 => x"58220018",
    15138 => x"58200010", 15139 => x"78010001", 15140 => x"38218f48",
    15141 => x"28210000", 15142 => x"28220000", 15143 => x"38420004",
    15144 => x"58220000", 15145 => x"34010000", 15146 => x"c3a00000",
    15147 => x"78050001", 15148 => x"38a58f48", 15149 => x"28a50000",
    15150 => x"202100ff", 15151 => x"00630003", 15152 => x"58a20014",
    15153 => x"58a10018", 15154 => x"58a30010", 15155 => x"34010003",
    15156 => x"5c810007", 15157 => x"28a20000", 15158 => x"3401fff3",
    15159 => x"a0410800", 15160 => x"38210008", 15161 => x"58a10000",
    15162 => x"c3a00000", 15163 => x"34010001", 15164 => x"5c810007",
    15165 => x"28a2001c", 15166 => x"3401ffe7", 15167 => x"a0410800",
    15168 => x"38210008", 15169 => x"58a1001c", 15170 => x"c3a00000",
    15171 => x"34010002", 15172 => x"5c810006", 15173 => x"28a2001c",
    15174 => x"3401ffe7", 15175 => x"a0410800", 15176 => x"38210010",
    15177 => x"58a1001c", 15178 => x"c3a00000", 15179 => x"379cffe0",
    15180 => x"5b8b0020", 15181 => x"5b8c001c", 15182 => x"5b8d0018",
    15183 => x"5b8e0014", 15184 => x"5b8f0010", 15185 => x"5b90000c",
    15186 => x"5b910008", 15187 => x"5b9d0004", 15188 => x"b8206000",
    15189 => x"78010001", 15190 => x"38215a88", 15191 => x"282f0000",
    15192 => x"780b0001", 15193 => x"b8406800", 15194 => x"396b8f48",
    15195 => x"fbffff9a", 15196 => x"b8208800", 15197 => x"29610000",
    15198 => x"b8408000", 15199 => x"282e0004", 15200 => x"a1cf7000",
    15201 => x"fbffff94", 15202 => x"5c31fff9", 15203 => x"5c50fff8",
    15204 => x"45800003", 15205 => x"59810000", 15206 => x"59820004",
    15207 => x"45a00003", 15208 => x"3dc10003", 15209 => x"59a10000",
    15210 => x"2b9d0004", 15211 => x"2b8b0020", 15212 => x"2b8c001c",
    15213 => x"2b8d0018", 15214 => x"2b8e0014", 15215 => x"2b8f0010",
    15216 => x"2b90000c", 15217 => x"2b910008", 15218 => x"379c0020",
    15219 => x"c3a00000", 15220 => x"78010001", 15221 => x"38218f48",
    15222 => x"28210000", 15223 => x"28210000", 15224 => x"20210004",
    15225 => x"64210000", 15226 => x"c3a00000", 15227 => x"78020001",
    15228 => x"38428f48", 15229 => x"28420000", 15230 => x"2843001c",
    15231 => x"44200003", 15232 => x"38630006", 15233 => x"e0000003",
    15234 => x"3401fff9", 15235 => x"a0611800", 15236 => x"5843001c",
    15237 => x"34010000", 15238 => x"c3a00000", 15239 => x"379cffe0",
    15240 => x"5b8b001c", 15241 => x"5b8c0018", 15242 => x"5b8d0014",
    15243 => x"5b8e0010", 15244 => x"5b8f000c", 15245 => x"5b900008",
    15246 => x"5b9d0004", 15247 => x"b8205800", 15248 => x"78010001",
    15249 => x"38218efc", 15250 => x"b8406000", 15251 => x"40220000",
    15252 => x"b8607000", 15253 => x"b8807800", 15254 => x"b8a06800",
    15255 => x"3401ffff", 15256 => x"4440002b", 15257 => x"3d8c0001",
    15258 => x"b9600800", 15259 => x"fbfff91b", 15260 => x"218200fe",
    15261 => x"b9600800", 15262 => x"fbfff960", 15263 => x"01c20008",
    15264 => x"b9600800", 15265 => x"204200ff", 15266 => x"fbfff95c",
    15267 => x"21c200ff", 15268 => x"b9600800", 15269 => x"fbfff959",
    15270 => x"b9600800", 15271 => x"fbfff923", 15272 => x"39820001",
    15273 => x"b9600800", 15274 => x"204200ff", 15275 => x"fbfff953",
    15276 => x"340c0000", 15277 => x"35aeffff", 15278 => x"37900023",
    15279 => x"e0000009", 15280 => x"b9600800", 15281 => x"ba001000",
    15282 => x"34030000", 15283 => x"fbfff988", 15284 => x"43820023",
    15285 => x"b5ec0800", 15286 => x"358c0001", 15287 => x"30220000",
    15288 => x"55ccfff8", 15289 => x"b9600800", 15290 => x"ba001000",
    15291 => x"34030001", 15292 => x"fbfff97f", 15293 => x"43810023",
    15294 => x"b5ee7000", 15295 => x"31c10000", 15296 => x"b9600800",
    15297 => x"fbfff925", 15298 => x"b9a00800", 15299 => x"2b9d0004",
    15300 => x"2b8b001c", 15301 => x"2b8c0018", 15302 => x"2b8d0014",
    15303 => x"2b8e0010", 15304 => x"2b8f000c", 15305 => x"2b900008",
    15306 => x"379c0020", 15307 => x"c3a00000", 15308 => x"379cffe0",
    15309 => x"5b8b0020", 15310 => x"5b8c001c", 15311 => x"5b8d0018",
    15312 => x"5b8e0014", 15313 => x"5b8f0010", 15314 => x"5b90000c",
    15315 => x"5b910008", 15316 => x"5b9d0004", 15317 => x"b8205800",
    15318 => x"78010001", 15319 => x"38218efc", 15320 => x"b8606800",
    15321 => x"40230000", 15322 => x"3c4f0001", 15323 => x"b8808000",
    15324 => x"b8a07000", 15325 => x"3401ffff", 15326 => x"21ef00ff",
    15327 => x"340c0000", 15328 => x"5c60001f", 15329 => x"e0000020",
    15330 => x"b9600800", 15331 => x"fbfff8d3", 15332 => x"b9e01000",
    15333 => x"b9600800", 15334 => x"fbfff918", 15335 => x"01a20008",
    15336 => x"b9600800", 15337 => x"204200ff", 15338 => x"fbfff914",
    15339 => x"21a200ff", 15340 => x"b9600800", 15341 => x"fbfff911",
    15342 => x"b60c1000", 15343 => x"40420000", 15344 => x"b9600800",
    15345 => x"35ad0001", 15346 => x"fbfff90c", 15347 => x"b9600800",
    15348 => x"fbfff8f2", 15349 => x"b9600800", 15350 => x"fbfff8c0",
    15351 => x"b9600800", 15352 => x"b9e01000", 15353 => x"fbfff905",
    15354 => x"b8208800", 15355 => x"b9600800", 15356 => x"fbfff8ea",
    15357 => x"5e20fff8", 15358 => x"358c0001", 15359 => x"55ccffe3",
    15360 => x"b9c00800", 15361 => x"2b9d0004", 15362 => x"2b8b0020",
    15363 => x"2b8c001c", 15364 => x"2b8d0018", 15365 => x"2b8e0014",
    15366 => x"2b8f0010", 15367 => x"2b90000c", 15368 => x"2b910008",
    15369 => x"379c0020", 15370 => x"c3a00000", 15371 => x"379cffec",
    15372 => x"5b8b0014", 15373 => x"5b8c0010", 15374 => x"5b8d000c",
    15375 => x"5b8e0008", 15376 => x"5b9d0004", 15377 => x"780d0001",
    15378 => x"780c0001", 15379 => x"39ad8f00", 15380 => x"398c8f04",
    15381 => x"780b0001", 15382 => x"59a10000", 15383 => x"59820000",
    15384 => x"34030001", 15385 => x"396b8efc", 15386 => x"202100ff",
    15387 => x"204200ff", 15388 => x"31630000", 15389 => x"fbfff97c",
    15390 => x"b8207000", 15391 => x"5c200006", 15392 => x"41a10003",
    15393 => x"41820003", 15394 => x"fbfff977", 15395 => x"5c2e0002",
    15396 => x"31600000", 15397 => x"2b9d0004", 15398 => x"2b8b0014",
    15399 => x"2b8c0010", 15400 => x"2b8d000c", 15401 => x"2b8e0008",
    15402 => x"379c0014", 15403 => x"c3a00000", 15404 => x"379cfff8",
    15405 => x"5b8b0008", 15406 => x"5b9d0004", 15407 => x"78010001",
    15408 => x"78020001", 15409 => x"38218f00", 15410 => x"38428f04",
    15411 => x"40420003", 15412 => x"780b0001", 15413 => x"40210003",
    15414 => x"396b71a8", 15415 => x"34031004", 15416 => x"b9602000",
    15417 => x"34050001", 15418 => x"31600000", 15419 => x"fbffff91",
    15420 => x"34030001", 15421 => x"3402ffff", 15422 => x"5c230002",
    15423 => x"41620000", 15424 => x"b8400800", 15425 => x"2b9d0004",
    15426 => x"2b8b0008", 15427 => x"379c0008", 15428 => x"c3a00000",
    15429 => x"379cffc4", 15430 => x"5b8b001c", 15431 => x"5b8c0018",
    15432 => x"5b8d0014", 15433 => x"5b8e0010", 15434 => x"5b8f000c",
    15435 => x"5b900008", 15436 => x"5b9d0004", 15437 => x"b8205800",
    15438 => x"206d00ff", 15439 => x"34010002", 15440 => x"204c00ff",
    15441 => x"3405fffc", 15442 => x"55a10087", 15443 => x"78040001",
    15444 => x"388471a8", 15445 => x"40820000", 15446 => x"340100ff",
    15447 => x"5c41000d", 15448 => x"78010001", 15449 => x"78020001",
    15450 => x"38218f00", 15451 => x"38428f04", 15452 => x"40420003",
    15453 => x"40210003", 15454 => x"34050001", 15455 => x"34031004",
    15456 => x"fbffff27", 15457 => x"34020001", 15458 => x"3405ffff",
    15459 => x"5c220076", 15460 => x"78010001", 15461 => x"382171a8",
    15462 => x"40230000", 15463 => x"340200ff", 15464 => x"5c620002",
    15465 => x"30200000", 15466 => x"5d800021", 15467 => x"78010001",
    15468 => x"382171a8", 15469 => x"40210000", 15470 => x"34050000",
    15471 => x"442c006a", 15472 => x"78010001", 15473 => x"78020001",
    15474 => x"38218f00", 15475 => x"38428f04", 15476 => x"09a3001d",
    15477 => x"40420003", 15478 => x"40210003", 15479 => x"3405001d",
    15480 => x"34631005", 15481 => x"b9602000", 15482 => x"fbffff0d",
    15483 => x"3402001d", 15484 => x"b9606000", 15485 => x"3405ffff",
    15486 => x"5c22005b", 15487 => x"3562001c", 15488 => x"34010000",
    15489 => x"e0000005", 15490 => x"41830000", 15491 => x"358c0001",
    15492 => x"b4230800", 15493 => x"202100ff", 15494 => x"5d82fffc",
    15495 => x"4162001c", 15496 => x"3405fffd", 15497 => x"5c410050",
    15498 => x"e000004a", 15499 => x"34010001", 15500 => x"5d810048",
    15501 => x"780f0001", 15502 => x"780e0001", 15503 => x"780d0001",
    15504 => x"340c0000", 15505 => x"39ef71a8", 15506 => x"39ce8f00",
    15507 => x"39ad8f04", 15508 => x"37900020", 15509 => x"e0000015",
    15510 => x"0983001d", 15511 => x"41a20003", 15512 => x"41c10003",
    15513 => x"34631005", 15514 => x"ba002000", 15515 => x"3405001d",
    15516 => x"fbfffeeb", 15517 => x"3402001d", 15518 => x"5c22003a",
    15519 => x"ba000800", 15520 => x"b9601000", 15521 => x"34030010",
    15522 => x"f8001084", 15523 => x"5c200005", 15524 => x"78010001",
    15525 => x"38215838", 15526 => x"fbfff549", 15527 => x"e0000005",
    15528 => x"358c0001", 15529 => x"218c00ff", 15530 => x"41e10000",
    15531 => x"542cffeb", 15532 => x"34010002", 15533 => x"3405fffe",
    15534 => x"5581002b", 15535 => x"3563001c", 15536 => x"b9600800",
    15537 => x"34020000", 15538 => x"e0000005", 15539 => x"40240000",
    15540 => x"34210001", 15541 => x"b4441000", 15542 => x"204200ff",
    15543 => x"5c23fffc", 15544 => x"780e0001", 15545 => x"780d0001",
    15546 => x"3162001c", 15547 => x"39ce8f00", 15548 => x"39ad8f04",
    15549 => x"0983001d", 15550 => x"41c10003", 15551 => x"41a20003",
    15552 => x"b9602000", 15553 => x"34631005", 15554 => x"3405001d",
    15555 => x"780b0001", 15556 => x"fbffff08", 15557 => x"396b71a8",
    15558 => x"41610000", 15559 => x"542c000d", 15560 => x"78010001",
    15561 => x"38215854", 15562 => x"fbfff525", 15563 => x"41610000",
    15564 => x"41a20003", 15565 => x"34031004", 15566 => x"34210001",
    15567 => x"31610000", 15568 => x"41c10003", 15569 => x"b9602000",
    15570 => x"34050001", 15571 => x"fbfffef9", 15572 => x"78010001",
    15573 => x"382171a8", 15574 => x"40250000", 15575 => x"e0000002",
    15576 => x"3405ffff", 15577 => x"b8a00800", 15578 => x"2b9d0004",
    15579 => x"2b8b001c", 15580 => x"2b8c0018", 15581 => x"2b8d0014",
    15582 => x"2b8e0010", 15583 => x"2b8f000c", 15584 => x"2b900008",
    15585 => x"379c003c", 15586 => x"c3a00000", 15587 => x"379cffcc",
    15588 => x"5b8b0014", 15589 => x"5b8c0010", 15590 => x"5b8d000c",
    15591 => x"5b8e0008", 15592 => x"5b9d0004", 15593 => x"340d0000",
    15594 => x"b8205800", 15595 => x"340c0001", 15596 => x"378e0018",
    15597 => x"e0000027", 15598 => x"b9c00800", 15599 => x"34020000",
    15600 => x"b9a01800", 15601 => x"fbffff54", 15602 => x"b8206000",
    15603 => x"4c010023", 15604 => x"b9c00800", 15605 => x"b9601000",
    15606 => x"34030010", 15607 => x"f800102f", 15608 => x"35ad0001",
    15609 => x"5c20001b", 15610 => x"2b81002c", 15611 => x"340c0001",
    15612 => x"00220018", 15613 => x"31610017", 15614 => x"31620014",
    15615 => x"00220010", 15616 => x"31620015", 15617 => x"00220008",
    15618 => x"2b810030", 15619 => x"31620016", 15620 => x"00220018",
    15621 => x"3161001b", 15622 => x"31620018", 15623 => x"00220010",
    15624 => x"31620019", 15625 => x"00220008", 15626 => x"2b810028",
    15627 => x"3162001a", 15628 => x"00220018", 15629 => x"31610013",
    15630 => x"31620010", 15631 => x"00220010", 15632 => x"31620011",
    15633 => x"00220008", 15634 => x"31620012", 15635 => x"e0000003",
    15636 => x"498dffda", 15637 => x"340c0000", 15638 => x"b9800800",
    15639 => x"2b9d0004", 15640 => x"2b8b0014", 15641 => x"2b8c0010",
    15642 => x"2b8d000c", 15643 => x"2b8e0008", 15644 => x"379c0034",
    15645 => x"c3a00000", 15646 => x"379cfff8", 15647 => x"5b8b0008",
    15648 => x"5b9d0004", 15649 => x"78030001", 15650 => x"b8205800",
    15651 => x"204200ff", 15652 => x"78010001", 15653 => x"38218f00",
    15654 => x"38638f04", 15655 => x"44400015", 15656 => x"29640000",
    15657 => x"78028000", 15658 => x"34050004", 15659 => x"b8821000",
    15660 => x"59620000", 15661 => x"40620003", 15662 => x"40210003",
    15663 => x"34031000", 15664 => x"b9602000", 15665 => x"fbfffe9b",
    15666 => x"7c210004", 15667 => x"78040001", 15668 => x"38845a68",
    15669 => x"c8011000", 15670 => x"29630000", 15671 => x"28810000",
    15672 => x"38420001", 15673 => x"a0610800", 15674 => x"59610000",
    15675 => x"e0000013", 15676 => x"40620003", 15677 => x"40210003",
    15678 => x"34031000", 15679 => x"b9602000", 15680 => x"34050004",
    15681 => x"fbfffe46", 15682 => x"34030004", 15683 => x"3402ffff",
    15684 => x"5c23000a", 15685 => x"29610000", 15686 => x"34020000",
    15687 => x"4c200007", 15688 => x"78030001", 15689 => x"38635a68",
    15690 => x"28620000", 15691 => x"a0220800", 15692 => x"59610000",
    15693 => x"34020001", 15694 => x"b8400800", 15695 => x"2b9d0004",
    15696 => x"2b8b0008", 15697 => x"379c0008", 15698 => x"c3a00000",
    15699 => x"379cfff8", 15700 => x"5b9d0004", 15701 => x"78010001",
    15702 => x"78020001", 15703 => x"38218f00", 15704 => x"38428f04",
    15705 => x"40420003", 15706 => x"40210003", 15707 => x"34031074",
    15708 => x"3784000a", 15709 => x"34050002", 15710 => x"0f80000a",
    15711 => x"fbfffe6d", 15712 => x"34030002", 15713 => x"3402ffff",
    15714 => x"5c230002", 15715 => x"2f82000a", 15716 => x"b8400800",
    15717 => x"2b9d0004", 15718 => x"379c0008", 15719 => x"c3a00000",
    15720 => x"379cffcc", 15721 => x"5b8b002c", 15722 => x"5b8c0028",
    15723 => x"5b8d0024", 15724 => x"5b8e0020", 15725 => x"5b8f001c",
    15726 => x"5b900018", 15727 => x"5b910014", 15728 => x"5b920010",
    15729 => x"5b93000c", 15730 => x"5b940008", 15731 => x"5b9d0004",
    15732 => x"78030001", 15733 => x"78020001", 15734 => x"38638f00",
    15735 => x"b8208800", 15736 => x"38428f04", 15737 => x"34010020",
    15738 => x"33810037", 15739 => x"40420003", 15740 => x"40610003",
    15741 => x"37840034", 15742 => x"34031074", 15743 => x"34050002",
    15744 => x"fbfffe07", 15745 => x"34020002", 15746 => x"340bffff",
    15747 => x"5c220051", 15748 => x"2f820034", 15749 => x"3801ffff",
    15750 => x"5c410002", 15751 => x"0f800034", 15752 => x"780d0001",
    15753 => x"780c0001", 15754 => x"340b0001", 15755 => x"39ad8f00",
    15756 => x"398c8f04", 15757 => x"37900037", 15758 => x"e0000023",
    15759 => x"41b40003", 15760 => x"41930003", 15761 => x"b9c00800",
    15762 => x"34721076", 15763 => x"f8000f64", 15764 => x"b8202800",
    15765 => x"b9c02000", 15766 => x"ba800800", 15767 => x"ba601000",
    15768 => x"ba401800", 15769 => x"fbfffe33", 15770 => x"b8207000",
    15771 => x"29e10000", 15772 => x"f8000f5b", 15773 => x"5dc10036",
    15774 => x"29e10000", 15775 => x"2f8e0034", 15776 => x"f8000f57",
    15777 => x"b5c11800", 15778 => x"41820003", 15779 => x"41a10003",
    15780 => x"2063ffff", 15781 => x"0f830034", 15782 => x"ba002000",
    15783 => x"34631076", 15784 => x"34050001", 15785 => x"fbfffe23",
    15786 => x"34020001", 15787 => x"5c220028", 15788 => x"2f810034",
    15789 => x"356b0001", 15790 => x"216b00ff", 15791 => x"34210001",
    15792 => x"0f810034", 15793 => x"3d6f0002", 15794 => x"2f830034",
    15795 => x"b62f7800", 15796 => x"29ee0000", 15797 => x"5dc0ffda",
    15798 => x"3401000a", 15799 => x"33810037", 15800 => x"41820003",
    15801 => x"41a10003", 15802 => x"34631075", 15803 => x"37840037",
    15804 => x"34050001", 15805 => x"fbfffe0f", 15806 => x"34020001",
    15807 => x"340bffff", 15808 => x"5c220014", 15809 => x"41a10003",
    15810 => x"41820003", 15811 => x"34031074", 15812 => x"37840034",
    15813 => x"34050002", 15814 => x"fbfffe06", 15815 => x"b8207000",
    15816 => x"34010002", 15817 => x"5dc1000b", 15818 => x"41a10003",
    15819 => x"41820003", 15820 => x"34031074", 15821 => x"37840032",
    15822 => x"34050002", 15823 => x"fbfffdb8", 15824 => x"e42e5800",
    15825 => x"356bffff", 15826 => x"e0000002", 15827 => x"340bffff",
    15828 => x"b9600800", 15829 => x"2b9d0004", 15830 => x"2b8b002c",
    15831 => x"2b8c0028", 15832 => x"2b8d0024", 15833 => x"2b8e0020",
    15834 => x"2b8f001c", 15835 => x"2b900018", 15836 => x"2b910014",
    15837 => x"2b920010", 15838 => x"2b93000c", 15839 => x"2b940008",
    15840 => x"379c0034", 15841 => x"c3a00000", 15842 => x"379cffe4",
    15843 => x"5b8b0018", 15844 => x"5b8c0014", 15845 => x"5b8d0010",
    15846 => x"5b8e000c", 15847 => x"5b8f0008", 15848 => x"5b9d0004",
    15849 => x"78010001", 15850 => x"78020001", 15851 => x"38218f00",
    15852 => x"38428f04", 15853 => x"40420003", 15854 => x"40210003",
    15855 => x"34031074", 15856 => x"3784001c", 15857 => x"34050002",
    15858 => x"fbfffd95", 15859 => x"34030002", 15860 => x"3402ffff",
    15861 => x"5c230025", 15862 => x"2f81001c", 15863 => x"3802fffd",
    15864 => x"3421ffff", 15865 => x"2021ffff", 15866 => x"50410005",
    15867 => x"78010001", 15868 => x"38214ec8", 15869 => x"0f80001c",
    15870 => x"fbfff3f1", 15871 => x"780e0001", 15872 => x"780d0001",
    15873 => x"780c0001", 15874 => x"340b0000", 15875 => x"39ce8f00",
    15876 => x"39ad8f04", 15877 => x"378f001f", 15878 => x"398c4ec4",
    15879 => x"e000000e", 15880 => x"41a20003", 15881 => x"41c10003",
    15882 => x"35631076", 15883 => x"b9e02000", 15884 => x"34050001",
    15885 => x"fbfffd7a", 15886 => x"34020001", 15887 => x"5c22000a",
    15888 => x"4382001f", 15889 => x"b9800800", 15890 => x"356b0001",
    15891 => x"fbfff3dc", 15892 => x"216bffff", 15893 => x"2f81001c",
    15894 => x"542bfff2", 15895 => x"34020000", 15896 => x"e0000002",
    15897 => x"3402ffff", 15898 => x"b8400800", 15899 => x"2b9d0004",
    15900 => x"2b8b0018", 15901 => x"2b8c0014", 15902 => x"2b8d0010",
    15903 => x"2b8e000c", 15904 => x"2b8f0008", 15905 => x"379c001c",
    15906 => x"c3a00000", 15907 => x"379cffdc", 15908 => x"5b8b0024",
    15909 => x"5b8c0020", 15910 => x"5b8d001c", 15911 => x"5b8e0018",
    15912 => x"5b8f0014", 15913 => x"5b900010", 15914 => x"5b91000c",
    15915 => x"5b920008", 15916 => x"5b9d0004", 15917 => x"206300ff",
    15918 => x"b8208800", 15919 => x"205200ff", 15920 => x"5c600012",
    15921 => x"78040001", 15922 => x"78030001", 15923 => x"38848f00",
    15924 => x"38638f04", 15925 => x"40620003", 15926 => x"40810003",
    15927 => x"78040001", 15928 => x"34031074", 15929 => x"38848f08",
    15930 => x"34050002", 15931 => x"fbfffd4c", 15932 => x"34020002",
    15933 => x"3403ffff", 15934 => x"5c22002b", 15935 => x"78030001",
    15936 => x"38638f0a", 15937 => x"0c610000", 15938 => x"78040001",
    15939 => x"38848f0a", 15940 => x"78030001", 15941 => x"38638f08",
    15942 => x"2c820000", 15943 => x"2c610000", 15944 => x"34030000",
    15945 => x"3442fffe", 15946 => x"5041001f", 15947 => x"780d0001",
    15948 => x"780c0001", 15949 => x"340b0000", 15950 => x"b8807000",
    15951 => x"39ad8f00", 15952 => x"398c8f04", 15953 => x"3410000a",
    15954 => x"2dc30000", 15955 => x"3461fffe", 15956 => x"54320012",
    15957 => x"41820003", 15958 => x"41a10003", 15959 => x"34640001",
    15960 => x"b62b7800", 15961 => x"0dc40000", 15962 => x"34631074",
    15963 => x"b9e02000", 15964 => x"34050001", 15965 => x"fbfffd2a",
    15966 => x"34020001", 15967 => x"5c220009", 15968 => x"41e10000",
    15969 => x"356b0001", 15970 => x"216b00ff", 15971 => x"5c30ffef",
    15972 => x"b9601800", 15973 => x"e0000004", 15974 => x"3403fffd",
    15975 => x"e0000002", 15976 => x"3403ffff", 15977 => x"b8600800",
    15978 => x"2b9d0004", 15979 => x"2b8b0024", 15980 => x"2b8c0020",
    15981 => x"2b8d001c", 15982 => x"2b8e0018", 15983 => x"2b8f0014",
    15984 => x"2b900010", 15985 => x"2b91000c", 15986 => x"2b920008",
    15987 => x"379c0024", 15988 => x"c3a00000", 15989 => x"379cfffc",
    15990 => x"5b9d0004", 15991 => x"78010001", 15992 => x"3821586c",
    15993 => x"fbfff376", 15994 => x"3401ffff", 15995 => x"2b9d0004",
    15996 => x"379c0004", 15997 => x"c3a00000", 15998 => x"379cfff8",
    15999 => x"5b8b0008", 16000 => x"5b9d0004", 16001 => x"78010001",
    16002 => x"b8405800", 16003 => x"78020001", 16004 => x"38425e48",
    16005 => x"38215890", 16006 => x"fbfff369", 16007 => x"78020001",
    16008 => x"78010001", 16009 => x"384291d0", 16010 => x"382191e0",
    16011 => x"34460090", 16012 => x"34050022", 16013 => x"34040033",
    16014 => x"28220004", 16015 => x"204300ff", 16016 => x"7c670042",
    16017 => x"7c630028", 16018 => x"a0e31800", 16019 => x"5c60000b",
    16020 => x"28230000", 16021 => x"31650000", 16022 => x"31640001",
    16023 => x"31630002", 16024 => x"00430018", 16025 => x"31630003",
    16026 => x"00430010", 16027 => x"00420008", 16028 => x"31630004",
    16029 => x"31620005", 16030 => x"34210010", 16031 => x"5c26ffef",
    16032 => x"34010000", 16033 => x"2b9d0004", 16034 => x"2b8b0008",
    16035 => x"379c0008", 16036 => x"c3a00000", 16037 => x"379cffe8",
    16038 => x"5b8b0018", 16039 => x"5b8c0014", 16040 => x"5b8d0010",
    16041 => x"5b8e000c", 16042 => x"5b8f0008", 16043 => x"5b9d0004",
    16044 => x"780b0001", 16045 => x"b8207800", 16046 => x"b8407000",
    16047 => x"340d0008", 16048 => x"340c0001", 16049 => x"396b71ac",
    16050 => x"a18e1800", 16051 => x"29640008", 16052 => x"7c620000",
    16053 => x"b9e00800", 16054 => x"35adffff", 16055 => x"d8800000",
    16056 => x"3d8c0001", 16057 => x"5da0fff9", 16058 => x"2b9d0004",
    16059 => x"2b8b0018", 16060 => x"2b8c0014", 16061 => x"2b8d0010",
    16062 => x"2b8e000c", 16063 => x"2b8f0008", 16064 => x"379c0018",
    16065 => x"c3a00000", 16066 => x"379cffe8", 16067 => x"5b8b0018",
    16068 => x"5b8c0014", 16069 => x"5b8d0010", 16070 => x"5b8e000c",
    16071 => x"5b8f0008", 16072 => x"5b9d0004", 16073 => x"780b0001",
    16074 => x"b8207800", 16075 => x"340e0008", 16076 => x"340c0000",
    16077 => x"340d0001", 16078 => x"396b71ac", 16079 => x"29620004",
    16080 => x"b9e00800", 16081 => x"35ceffff", 16082 => x"d8400000",
    16083 => x"7c220000", 16084 => x"c8021000", 16085 => x"a1a21000",
    16086 => x"b9826000", 16087 => x"3dad0001", 16088 => x"5dc0fff7",
    16089 => x"34010064", 16090 => x"fbffe980", 16091 => x"b9800800",
    16092 => x"2b9d0004", 16093 => x"2b8b0018", 16094 => x"2b8c0014",
    16095 => x"2b8d0010", 16096 => x"2b8e000c", 16097 => x"2b8f0008",
    16098 => x"379c0018", 16099 => x"c3a00000", 16100 => x"379cffc0",
    16101 => x"5b8b0040", 16102 => x"5b8c003c", 16103 => x"5b8d0038",
    16104 => x"5b8e0034", 16105 => x"5b8f0030", 16106 => x"5b90002c",
    16107 => x"5b910028", 16108 => x"5b920024", 16109 => x"5b930020",
    16110 => x"5b94001c", 16111 => x"5b950018", 16112 => x"5b960014",
    16113 => x"5b970010", 16114 => x"5b98000c", 16115 => x"5b990008",
    16116 => x"5b9d0004", 16117 => x"34020000", 16118 => x"b8206000",
    16119 => x"34030080", 16120 => x"34210008", 16121 => x"780d0001",
    16122 => x"f8000d47", 16123 => x"39ad71ac", 16124 => x"29a10000",
    16125 => x"340f0000", 16126 => x"44200061", 16127 => x"b9805800",
    16128 => x"34120000", 16129 => x"34110000", 16130 => x"78194000",
    16131 => x"34160001", 16132 => x"34180008", 16133 => x"596c0008",
    16134 => x"45e00022", 16135 => x"29610000", 16136 => x"78028000",
    16137 => x"34030000", 16138 => x"59610010", 16139 => x"29610004",
    16140 => x"59610014", 16141 => x"a0590800", 16142 => x"44200003",
    16143 => x"78024000", 16144 => x"34030000", 16145 => x"a0710800",
    16146 => x"a0522800", 16147 => x"b8a12800", 16148 => x"29640010",
    16149 => x"29610014", 16150 => x"5ca0000e", 16151 => x"a4603000",
    16152 => x"a0260800", 16153 => x"59610014", 16154 => x"00630001",
    16155 => x"3c41001f", 16156 => x"a4403800", 16157 => x"00420001",
    16158 => x"a0872000", 16159 => x"b8231800", 16160 => x"59640010",
    16161 => x"b8430800", 16162 => x"5c25ffeb", 16163 => x"e000003c",
    16164 => x"b8821000", 16165 => x"b8231800", 16166 => x"59620010",
    16167 => x"59630014", 16168 => x"35ee0001", 16169 => x"29a20000",
    16170 => x"3dce0004", 16171 => x"b9800800", 16172 => x"b58e7000",
    16173 => x"d8400000", 16174 => x"5c360031", 16175 => x"b9800800",
    16176 => x"340200f0", 16177 => x"fbffff74", 16178 => x"34140040",
    16179 => x"34130000", 16180 => x"34100001", 16181 => x"34120000",
    16182 => x"34110000", 16183 => x"29a20004", 16184 => x"b9800800",
    16185 => x"29d70004", 16186 => x"d8400000", 16187 => x"29a20004",
    16188 => x"b820a800", 16189 => x"b9800800", 16190 => x"a2f0b800",
    16191 => x"d8400000", 16192 => x"46a10008", 16193 => x"29a30008",
    16194 => x"baa01000", 16195 => x"7eb50000", 16196 => x"b9800800",
    16197 => x"d8600000", 16198 => x"5eb60011", 16199 => x"e0000007",
    16200 => x"29a30008", 16201 => x"b9800800", 16202 => x"bae01000",
    16203 => x"d8600000", 16204 => x"46e00009", 16205 => x"e000000a",
    16206 => x"29c10000", 16207 => x"b8330800", 16208 => x"59c10000",
    16209 => x"29c10004", 16210 => x"b8300800", 16211 => x"59c10004",
    16212 => x"e0000003", 16213 => x"ba539000", 16214 => x"ba308800",
    16215 => x"3e010001", 16216 => x"3e730001", 16217 => x"f6018000",
    16218 => x"3694ffff", 16219 => x"b6139800", 16220 => x"b8208000",
    16221 => x"5e80ffda", 16222 => x"e0000014", 16223 => x"b9e00800",
    16224 => x"2b9d0004", 16225 => x"2b8b0040", 16226 => x"2b8c003c",
    16227 => x"2b8d0038", 16228 => x"2b8e0034", 16229 => x"2b8f0030",
    16230 => x"2b90002c", 16231 => x"2b910028", 16232 => x"2b920024",
    16233 => x"2b930020", 16234 => x"2b94001c", 16235 => x"2b950018",
    16236 => x"2b960014", 16237 => x"2b970010", 16238 => x"2b98000c",
    16239 => x"2b990008", 16240 => x"379c0040", 16241 => x"c3a00000",
    16242 => x"35ef0001", 16243 => x"356b0010", 16244 => x"5df8ff91",
    16245 => x"e3ffffea", 16246 => x"379cfff0", 16247 => x"5b8b0010",
    16248 => x"5b8c000c", 16249 => x"5b8d0008", 16250 => x"5b9d0004",
    16251 => x"b8205800", 16252 => x"78010001", 16253 => x"382171ac",
    16254 => x"28220000", 16255 => x"29610000", 16256 => x"340c0000",
    16257 => x"340d0040", 16258 => x"d8400000", 16259 => x"29610000",
    16260 => x"34020055", 16261 => x"fbffff20", 16262 => x"29610008",
    16263 => x"2962000c", 16264 => x"b9801800", 16265 => x"358c0008",
    16266 => x"f8000b7c", 16267 => x"29610000", 16268 => x"fbffff19",
    16269 => x"5d8dfff9", 16270 => x"2b9d0004", 16271 => x"2b8b0010",
    16272 => x"2b8c000c", 16273 => x"2b8d0008", 16274 => x"379c0010",
    16275 => x"c3a00000", 16276 => x"28210000", 16277 => x"78020001",
    16278 => x"38429258", 16279 => x"28420000", 16280 => x"3c210008",
    16281 => x"3821000a", 16282 => x"58410000", 16283 => x"28410000",
    16284 => x"20230008", 16285 => x"5c60fffe", 16286 => x"20210001",
    16287 => x"18210001", 16288 => x"c3a00000", 16289 => x"28210000",
    16290 => x"78020001", 16291 => x"38429258", 16292 => x"28420000",
    16293 => x"3c210008", 16294 => x"38210009", 16295 => x"58410000",
    16296 => x"28410000", 16297 => x"20230008", 16298 => x"5c60fffe",
    16299 => x"20210001", 16300 => x"c3a00000", 16301 => x"28210000",
    16302 => x"78030001", 16303 => x"38639258", 16304 => x"3c210008",
    16305 => x"28630000", 16306 => x"7c420000", 16307 => x"38210008",
    16308 => x"b8221000", 16309 => x"58620000", 16310 => x"28610000",
    16311 => x"20210008", 16312 => x"5c20fffe", 16313 => x"c3a00000",
    16314 => x"78010001", 16315 => x"78030001", 16316 => x"38219258",
    16317 => x"38635aa4", 16318 => x"28210000", 16319 => x"28620000",
    16320 => x"58220004", 16321 => x"c3a00000", 16322 => x"379cffc4",
    16323 => x"5b8b001c", 16324 => x"5b8c0018", 16325 => x"5b8d0014",
    16326 => x"5b8e0010", 16327 => x"5b8f000c", 16328 => x"5b900008",
    16329 => x"5b9d0004", 16330 => x"b8206000", 16331 => x"28210000",
    16332 => x"340bffff", 16333 => x"4420002a", 16334 => x"29820004",
    16335 => x"44400028", 16336 => x"fbffe83e", 16337 => x"780e0001",
    16338 => x"b8206800", 16339 => x"340b0000", 16340 => x"3410001f",
    16341 => x"378f0020", 16342 => x"39ce58ac", 16343 => x"e000000b",
    16344 => x"fbffe836", 16345 => x"202400ff", 16346 => x"b56d1000",
    16347 => x"b5eb0800", 16348 => x"30240000", 16349 => x"b8401800",
    16350 => x"b9c00800", 16351 => x"b8802800", 16352 => x"fbfff20f",
    16353 => x"356b0001", 16354 => x"29810004", 16355 => x"ee0b1800",
    16356 => x"358c0004", 16357 => x"7c220000", 16358 => x"a0621000",
    16359 => x"5c40fff1", 16360 => x"78010001", 16361 => x"b9602000",
    16362 => x"b9a01000", 16363 => x"b9e01800", 16364 => x"382191d0",
    16365 => x"f80001cc", 16366 => x"b8206000", 16367 => x"b9601800",
    16368 => x"78010001", 16369 => x"fd8b5800", 16370 => x"382158d0",
    16371 => x"b9a01000", 16372 => x"b9802000", 16373 => x"fbfff1fa",
    16374 => x"c80b5800", 16375 => x"b9600800", 16376 => x"2b9d0004",
    16377 => x"2b8b001c", 16378 => x"2b8c0018", 16379 => x"2b8d0014",
    16380 => x"2b8e0010", 16381 => x"2b8f000c", 16382 => x"2b900008",
    16383 => x"379c003c", 16384 => x"c3a00000", 16385 => x"379cffc8",
    16386 => x"5b8b0018", 16387 => x"5b8c0014", 16388 => x"5b8d0010",
    16389 => x"5b8e000c", 16390 => x"5b8f0008", 16391 => x"5b9d0004",
    16392 => x"b8205800", 16393 => x"28210000", 16394 => x"3405ffff",
    16395 => x"4420002c", 16396 => x"29620004", 16397 => x"4440002a",
    16398 => x"fbffe800", 16399 => x"b8207000", 16400 => x"29610004",
    16401 => x"fbffe7fd", 16402 => x"b8205800", 16403 => x"34010020",
    16404 => x"4c2b0002", 16405 => x"340b0020", 16406 => x"378d001c",
    16407 => x"78010001", 16408 => x"b9602000", 16409 => x"b9c01000",
    16410 => x"b9a01800", 16411 => x"382191d0", 16412 => x"f8000189",
    16413 => x"b8206000", 16414 => x"78010001", 16415 => x"b9601800",
    16416 => x"382158f0", 16417 => x"b9c01000", 16418 => x"b9802000",
    16419 => x"fbfff1cc", 16420 => x"e98b5800", 16421 => x"ec0c0800",
    16422 => x"3405ffff", 16423 => x"b9615800", 16424 => x"5d60000f",
    16425 => x"b9a07800", 16426 => x"780d0001", 16427 => x"39ad58ac",
    16428 => x"b5eb0800", 16429 => x"40240000", 16430 => x"b56e1000",
    16431 => x"b9a00800", 16432 => x"b8401800", 16433 => x"b8802800",
    16434 => x"356b0001", 16435 => x"fbfff1bc", 16436 => x"498bfff8",
    16437 => x"fd8b2800", 16438 => x"c8052800", 16439 => x"b8a00800",
    16440 => x"2b9d0004", 16441 => x"2b8b0018", 16442 => x"2b8c0014",
    16443 => x"2b8d0010", 16444 => x"2b8e000c", 16445 => x"2b8f0008",
    16446 => x"379c0038", 16447 => x"c3a00000", 16448 => x"379cffe4",
    16449 => x"5b8b001c", 16450 => x"5b8c0018", 16451 => x"5b8d0014",
    16452 => x"5b8e0010", 16453 => x"5b8f000c", 16454 => x"5b900008",
    16455 => x"5b9d0004", 16456 => x"780d0001", 16457 => x"39ad91d0",
    16458 => x"b9a00800", 16459 => x"780b0001", 16460 => x"780f0001",
    16461 => x"780e0001", 16462 => x"fbfffe96", 16463 => x"396b91e0",
    16464 => x"340c0000", 16465 => x"39ef5910", 16466 => x"39ce5928",
    16467 => x"34100008", 16468 => x"29630000", 16469 => x"29640004",
    16470 => x"b8640800", 16471 => x"44200010", 16472 => x"b9801000",
    16473 => x"b9e00800", 16474 => x"fbfff195", 16475 => x"3d810004",
    16476 => x"34020000", 16477 => x"34210008", 16478 => x"b5a10800",
    16479 => x"f8000015", 16480 => x"2023ffff", 16481 => x"08632710",
    16482 => x"b8201000", 16483 => x"14420010", 16484 => x"14630010",
    16485 => x"b9c00800", 16486 => x"fbfff189", 16487 => x"358c0001",
    16488 => x"356b0010", 16489 => x"5d90ffeb", 16490 => x"34010000",
    16491 => x"2b9d0004", 16492 => x"2b8b001c", 16493 => x"2b8c0018",
    16494 => x"2b8d0014", 16495 => x"2b8e0010", 16496 => x"2b8f000c",
    16497 => x"2b900008", 16498 => x"379c001c", 16499 => x"c3a00000",
    16500 => x"379cffec", 16501 => x"5b8b0014", 16502 => x"5b8c0010",
    16503 => x"5b8d000c", 16504 => x"5b8e0008", 16505 => x"5b9d0004",
    16506 => x"402d000f", 16507 => x"b8206000", 16508 => x"34010028",
    16509 => x"b8407000", 16510 => x"45a10005", 16511 => x"34010042",
    16512 => x"45a10003", 16513 => x"34010010", 16514 => x"5da10034",
    16515 => x"21cb0002", 16516 => x"5d60000f", 16517 => x"b9800800",
    16518 => x"fbfffef0", 16519 => x"29810000", 16520 => x"34020044",
    16521 => x"21ce0001", 16522 => x"fbfffe1b", 16523 => x"34010000",
    16524 => x"5dcb002d", 16525 => x"780b0001", 16526 => x"396b71ac",
    16527 => x"29620004", 16528 => x"29810000", 16529 => x"d8400000",
    16530 => x"4420fffd", 16531 => x"b9800800", 16532 => x"fbfffee2",
    16533 => x"29810000", 16534 => x"780b0001", 16535 => x"340200be",
    16536 => x"396b8f0c", 16537 => x"fbfffe0c", 16538 => x"356e0008",
    16539 => x"e0000005", 16540 => x"29810000", 16541 => x"fbfffe25",
    16542 => x"31610000", 16543 => x"356b0001", 16544 => x"5d6efffc",
    16545 => x"78020001", 16546 => x"38428f0c", 16547 => x"40410001",
    16548 => x"40430000", 16549 => x"3c210008", 16550 => x"b8230800",
    16551 => x"34030028", 16552 => x"dc200800", 16553 => x"45a3000b",
    16554 => x"34030042", 16555 => x"45a30009", 16556 => x"34030010",
    16557 => x"5da3000b", 16558 => x"40420006", 16559 => x"3c21000f",
    16560 => x"3c42000c", 16561 => x"3421c000", 16562 => x"b8220800",
    16563 => x"e0000006", 16564 => x"3c21000c", 16565 => x"e0000004",
    16566 => x"78018000", 16567 => x"e0000002", 16568 => x"34010000",
    16569 => x"2b9d0004", 16570 => x"2b8b0014", 16571 => x"2b8c0010",
    16572 => x"2b8d000c", 16573 => x"2b8e0008", 16574 => x"379c0014",
    16575 => x"c3a00000", 16576 => x"379cfffc", 16577 => x"5b9d0004",
    16578 => x"34030000", 16579 => x"b8202000", 16580 => x"34090028",
    16581 => x"34080042", 16582 => x"34070010", 16583 => x"34060008",
    16584 => x"40850017", 16585 => x"44a90003", 16586 => x"44a80002",
    16587 => x"5ca70006", 16588 => x"3c630004", 16589 => x"34630008",
    16590 => x"b4230800", 16591 => x"fbffffa5", 16592 => x"e0000005",
    16593 => x"34630001", 16594 => x"34840010", 16595 => x"5c66fff5",
    16596 => x"78018000", 16597 => x"2b9d0004", 16598 => x"379c0004",
    16599 => x"c3a00000", 16600 => x"379cffe0", 16601 => x"5b8b0020",
    16602 => x"5b8c001c", 16603 => x"5b8d0018", 16604 => x"5b8e0014",
    16605 => x"5b8f0010", 16606 => x"5b90000c", 16607 => x"5b910008",
    16608 => x"5b9d0004", 16609 => x"b8205800", 16610 => x"b8408800",
    16611 => x"b8608000", 16612 => x"b8806000", 16613 => x"fbfffe91",
    16614 => x"29610000", 16615 => x"3402000f", 16616 => x"222e00ff",
    16617 => x"fbfffdbc", 16618 => x"29610000", 16619 => x"b9c01000",
    16620 => x"2231ff00", 16621 => x"fbfffdb8", 16622 => x"16310008",
    16623 => x"29610000", 16624 => x"ba201000", 16625 => x"340d0000",
    16626 => x"fbfffdb3", 16627 => x"e0000006", 16628 => x"b60d1000",
    16629 => x"29610000", 16630 => x"40420000", 16631 => x"35ad0001",
    16632 => x"fbfffdad", 16633 => x"498dfffb", 16634 => x"b9600800",
    16635 => x"fbfffe7b", 16636 => x"29610000", 16637 => x"340200aa",
    16638 => x"fbfffda7", 16639 => x"29610000", 16640 => x"fbfffdc2",
    16641 => x"b8207800", 16642 => x"5c2e0022", 16643 => x"29610000",
    16644 => x"fbfffdbe", 16645 => x"b8207000", 16646 => x"5c310020",
    16647 => x"29610000", 16648 => x"340d0000", 16649 => x"fbfffdb9",
    16650 => x"b8208800", 16651 => x"e0000007", 16652 => x"29610000",
    16653 => x"fbfffdb5", 16654 => x"b60d1000", 16655 => x"40420000",
    16656 => x"5c220018", 16657 => x"35ad0001", 16658 => x"498dfffa",
    16659 => x"b9600800", 16660 => x"fbfffe62", 16661 => x"29610000",
    16662 => x"34020055", 16663 => x"fbfffd8e", 16664 => x"29610000",
    16665 => x"b9e01000", 16666 => x"fbfffd8b", 16667 => x"29610000",
    16668 => x"b9c01000", 16669 => x"fbfffd88", 16670 => x"29610000",
    16671 => x"ba201000", 16672 => x"fbfffd85", 16673 => x"34012710",
    16674 => x"fbffe738", 16675 => x"e0000006", 16676 => x"340cffff",
    16677 => x"e0000004", 16678 => x"340cfffe", 16679 => x"e0000002",
    16680 => x"340cfffd", 16681 => x"b9800800", 16682 => x"2b9d0004",
    16683 => x"2b8b0020", 16684 => x"2b8c001c", 16685 => x"2b8d0018",
    16686 => x"2b8e0014", 16687 => x"2b8f0010", 16688 => x"2b90000c",
    16689 => x"2b910008", 16690 => x"379c0020", 16691 => x"c3a00000",
    16692 => x"379cffe4", 16693 => x"5b8b001c", 16694 => x"5b8c0018",
    16695 => x"5b8d0014", 16696 => x"5b8e0010", 16697 => x"5b8f000c",
    16698 => x"5b900008", 16699 => x"5b9d0004", 16700 => x"b8208000",
    16701 => x"2041001f", 16702 => x"b8405800", 16703 => x"b8607000",
    16704 => x"b8806000", 16705 => x"340d0000", 16706 => x"44200030",
    16707 => x"3441ffff", 16708 => x"b4240800", 16709 => x"1422001f",
    16710 => x"b8807800", 16711 => x"0042001b", 16712 => x"b4410800",
    16713 => x"1562001f", 16714 => x"14210005", 16715 => x"0042001b",
    16716 => x"b44b1000", 16717 => x"14420005", 16718 => x"4422000c",
    16719 => x"78010001", 16720 => x"38215aa8", 16721 => x"28220000",
    16722 => x"a1621000", 16723 => x"4c400005", 16724 => x"3442ffff",
    16725 => x"3401ffe0", 16726 => x"b8411000", 16727 => x"34420001",
    16728 => x"340f0020", 16729 => x"c9e27800", 16730 => x"ba000800",
    16731 => x"b9601000", 16732 => x"b9c01800", 16733 => x"b9e02000",
    16734 => x"fbffff7a", 16735 => x"b8206800", 16736 => x"48010016",
    16737 => x"b5cf7000", 16738 => x"b56f5800", 16739 => x"c98f6000",
    16740 => x"e000000e", 16741 => x"b9802000", 16742 => x"4dec0002",
    16743 => x"34040020", 16744 => x"ba000800", 16745 => x"b9601000",
    16746 => x"b9c01800", 16747 => x"fbffff6d", 16748 => x"48010009",
    16749 => x"b5a16800", 16750 => x"35ce0020", 16751 => x"356b0020",
    16752 => x"358cffe0", 16753 => x"e0000002", 16754 => x"340f0020",
    16755 => x"4980fff2", 16756 => x"e0000002", 16757 => x"b8206800",
    16758 => x"b9a00800", 16759 => x"2b9d0004", 16760 => x"2b8b001c",
    16761 => x"2b8c0018", 16762 => x"2b8d0014", 16763 => x"2b8e0010",
    16764 => x"2b8f000c", 16765 => x"2b900008", 16766 => x"379c001c",
    16767 => x"c3a00000", 16768 => x"379cffec", 16769 => x"5b8b0014",
    16770 => x"5b8c0010", 16771 => x"5b8d000c", 16772 => x"5b8e0008",
    16773 => x"5b9d0004", 16774 => x"b8405800", 16775 => x"b8206000",
    16776 => x"b8607000", 16777 => x"b8806800", 16778 => x"fbfffdec",
    16779 => x"29810000", 16780 => x"340200f0", 16781 => x"fbfffd18",
    16782 => x"29810000", 16783 => x"216200ff", 16784 => x"fbfffd15",
    16785 => x"2162ff00", 16786 => x"29810000", 16787 => x"00420008",
    16788 => x"340b0000", 16789 => x"fbfffd10", 16790 => x"e0000006",
    16791 => x"29810000", 16792 => x"fbfffd2a", 16793 => x"b5cb1000",
    16794 => x"30410000", 16795 => x"356b0001", 16796 => x"49abfffb",
    16797 => x"b9a00800", 16798 => x"2b9d0004", 16799 => x"2b8b0014",
    16800 => x"2b8c0010", 16801 => x"2b8d000c", 16802 => x"2b8e0008",
    16803 => x"379c0014", 16804 => x"c3a00000", 16805 => x"379cfffc",
    16806 => x"5b9d0004", 16807 => x"34050000", 16808 => x"b8203000",
    16809 => x"34080043", 16810 => x"34070008", 16811 => x"40c90017",
    16812 => x"5d280006", 16813 => x"3ca50004", 16814 => x"34a50008",
    16815 => x"b4250800", 16816 => x"fbffffd0", 16817 => x"e0000005",
    16818 => x"34a50001", 16819 => x"34c60010", 16820 => x"5ca7fff7",
    16821 => x"3401ffff", 16822 => x"2b9d0004", 16823 => x"379c0004",
    16824 => x"c3a00000", 16825 => x"379cfffc", 16826 => x"5b9d0004",
    16827 => x"34050000", 16828 => x"b8203000", 16829 => x"34080043",
    16830 => x"34070008", 16831 => x"40c90017", 16832 => x"5d280006",
    16833 => x"3ca50004", 16834 => x"34a50008", 16835 => x"b4250800",
    16836 => x"fbffff70", 16837 => x"e0000005", 16838 => x"34a50001",
    16839 => x"34c60010", 16840 => x"5ca7fff7", 16841 => x"3401ffff",
    16842 => x"2b9d0004", 16843 => x"379c0004", 16844 => x"c3a00000",
    16845 => x"379cfff4", 16846 => x"5b8b000c", 16847 => x"5b8c0008",
    16848 => x"5b9d0004", 16849 => x"780b0001", 16850 => x"396b8f1c",
    16851 => x"29610000", 16852 => x"5c200009", 16853 => x"fbfff5da",
    16854 => x"78020001", 16855 => x"342103e8", 16856 => x"38428f14",
    16857 => x"58410000", 16858 => x"29610000", 16859 => x"34210001",
    16860 => x"59610000", 16861 => x"780b0001", 16862 => x"396b8f18",
    16863 => x"296c0000", 16864 => x"fbfff5cf", 16865 => x"78020001",
    16866 => x"38428f14", 16867 => x"28440000", 16868 => x"c8242800",
    16869 => x"34010000", 16870 => x"48050018", 16871 => x"21830001",
    16872 => x"78010001", 16873 => x"3c650002", 16874 => x"38215e5c",
    16875 => x"b4250800", 16876 => x"28210000", 16877 => x"b4242000",
    16878 => x"29610000", 16879 => x"58440000", 16880 => x"34020001",
    16881 => x"34210001", 16882 => x"59610000", 16883 => x"78010001",
    16884 => x"382191d0", 16885 => x"44620003", 16886 => x"fbfffeca",
    16887 => x"e0000006", 16888 => x"34020002", 16889 => x"fbfffec7",
    16890 => x"78020001", 16891 => x"384271b8", 16892 => x"58410004",
    16893 => x"34010001", 16894 => x"2b9d0004", 16895 => x"2b8b000c",
    16896 => x"2b8c0008", 16897 => x"379c000c", 16898 => x"c3a00000",
    16899 => x"78010001", 16900 => x"38219288", 16901 => x"28220000",
    16902 => x"78010001", 16903 => x"382192b4", 16904 => x"58220000",
    16905 => x"340103c6", 16906 => x"58410004", 16907 => x"c3a00000",
    16908 => x"c3a00000", 16909 => x"379cfff8", 16910 => x"5b8b0008",
    16911 => x"5b9d0004", 16912 => x"b8205800", 16913 => x"3401000a",
    16914 => x"5d610003", 16915 => x"3401000d", 16916 => x"fbfffff9",
    16917 => x"78020001", 16918 => x"384292b4", 16919 => x"28420000",
    16920 => x"28410000", 16921 => x"20210001", 16922 => x"5c20fffe",
    16923 => x"584b0008", 16924 => x"2b9d0004", 16925 => x"2b8b0008",
    16926 => x"379c0008", 16927 => x"c3a00000", 16928 => x"379cfff4",
    16929 => x"5b8b000c", 16930 => x"5b8c0008", 16931 => x"5b9d0004",
    16932 => x"b8206000", 16933 => x"b8205800", 16934 => x"e0000004",
    16935 => x"b8400800", 16936 => x"356b0001", 16937 => x"fbffffe4",
    16938 => x"41620000", 16939 => x"5c40fffc", 16940 => x"c96c0800",
    16941 => x"2b9d0004", 16942 => x"2b8b000c", 16943 => x"2b8c0008",
    16944 => x"379c000c", 16945 => x"c3a00000", 16946 => x"78010001",
    16947 => x"382192b4", 16948 => x"28220000", 16949 => x"3401ffff",
    16950 => x"28430000", 16951 => x"20630002", 16952 => x"44600003",
    16953 => x"2841000c", 16954 => x"202100ff", 16955 => x"c3a00000",
    16956 => x"28250008", 16957 => x"28240000", 16958 => x"28260004",
    16959 => x"b4451800", 16960 => x"88642000", 16961 => x"5822001c",
    16962 => x"88461000", 16963 => x"b4821000", 16964 => x"2824000c",
    16965 => x"1442000c", 16966 => x"b4442000", 16967 => x"28220014",
    16968 => x"4c820005", 16969 => x"28240010", 16970 => x"44800008",
    16971 => x"4ca3000b", 16972 => x"e0000006", 16973 => x"28220018",
    16974 => x"4c440006", 16975 => x"28240010", 16976 => x"44800002",
    16977 => x"4c650005", 16978 => x"58230008", 16979 => x"e0000003",
    16980 => x"58230008", 16981 => x"b8801000", 16982 => x"58220020",
    16983 => x"b8400800", 16984 => x"c3a00000", 16985 => x"2822000c",
    16986 => x"58200008", 16987 => x"58220020", 16988 => x"c3a00000",
    16989 => x"379cfff8", 16990 => x"5b8b0008", 16991 => x"5b9d0004",
    16992 => x"b8205800", 16993 => x"58200014", 16994 => x"b8400800",
    16995 => x"f800093b", 16996 => x"2963000c", 16997 => x"29620000",
    16998 => x"4823000b", 16999 => x"29610004", 17000 => x"4c410003",
    17001 => x"34420001", 17002 => x"59620000", 17003 => x"29620000",
    17004 => x"5c410011", 17005 => x"34010001", 17006 => x"59610014",
    17007 => x"59610010", 17008 => x"e000000e", 17009 => x"29610008",
    17010 => x"4c220003", 17011 => x"3442ffff", 17012 => x"59620000",
    17013 => x"29620000", 17014 => x"5c410007", 17015 => x"34010001",
    17016 => x"59610014", 17017 => x"59600000", 17018 => x"59600010",
    17019 => x"3401ffff", 17020 => x"e0000002", 17021 => x"29610010",
    17022 => x"2b9d0004", 17023 => x"2b8b0008", 17024 => x"379c0008",
    17025 => x"c3a00000", 17026 => x"58200010", 17027 => x"58200000",
    17028 => x"58200014", 17029 => x"c3a00000", 17030 => x"78030001",
    17031 => x"38639294", 17032 => x"28640000", 17033 => x"48810013",
    17034 => x"78030001", 17035 => x"38638f30", 17036 => x"c8240800",
    17037 => x"44400007", 17038 => x"28620000", 17039 => x"34040001",
    17040 => x"bc810800", 17041 => x"28430028", 17042 => x"b8230800",
    17043 => x"e0000007", 17044 => x"28620000", 17045 => x"34040001",
    17046 => x"bc810800", 17047 => x"28430028", 17048 => x"a4200800",
    17049 => x"a0230800", 17050 => x"58410028", 17051 => x"c3a00000",
    17052 => x"78030001", 17053 => x"38638f30", 17054 => x"44400007",
    17055 => x"28620000", 17056 => x"34040001", 17057 => x"bc810800",
    17058 => x"28430024", 17059 => x"b8230800", 17060 => x"e0000007",
    17061 => x"28620000", 17062 => x"34040001", 17063 => x"bc810800",
    17064 => x"28430024", 17065 => x"a4200800", 17066 => x"a0230800",
    17067 => x"58410024", 17068 => x"c3a00000", 17069 => x"379cfff0",
    17070 => x"5b8b0010", 17071 => x"5b8c000c", 17072 => x"5b8d0008",
    17073 => x"5b9d0004", 17074 => x"b8406800", 17075 => x"b8606000",
    17076 => x"34020000", 17077 => x"34030028", 17078 => x"b8205800",
    17079 => x"f800098a", 17080 => x"b9600800", 17081 => x"b9a01000",
    17082 => x"34030014", 17083 => x"f8000908", 17084 => x"596c0014",
    17085 => x"2b9d0004", 17086 => x"2b8b0010", 17087 => x"2b8c000c",
    17088 => x"2b8d0008", 17089 => x"379c0010", 17090 => x"c3a00000",
    17091 => x"b8201800", 17092 => x"e0000004", 17093 => x"28840000",
    17094 => x"34630008", 17095 => x"44820006", 17096 => x"28610004",
    17097 => x"b8602000", 17098 => x"5c20fffb", 17099 => x"78010001",
    17100 => x"38215944", 17101 => x"c3a00000", 17102 => x"78020001",
    17103 => x"38428f30", 17104 => x"28420000", 17105 => x"b8201800",
    17106 => x"34010000", 17107 => x"28440008", 17108 => x"20840002",
    17109 => x"4480000c", 17110 => x"34040002", 17111 => x"58440008",
    17112 => x"78060001", 17113 => x"28420010", 17114 => x"38c65aac",
    17115 => x"28c40000", 17116 => x"3445ff9b", 17117 => x"54a40004",
    17118 => x"08420064", 17119 => x"34010001", 17120 => x"58620000",
    17121 => x"c3a00000", 17122 => x"379cfff0", 17123 => x"5b8b0010",
    17124 => x"5b8c000c", 17125 => x"5b8d0008", 17126 => x"5b9d0004",
    17127 => x"780b0001", 17128 => x"b8206000", 17129 => x"78010001",
    17130 => x"396b9294", 17131 => x"3821928c", 17132 => x"28210000",
    17133 => x"296d0000", 17134 => x"b42d6800", 17135 => x"29810000",
    17136 => x"b9a01000", 17137 => x"f8000114", 17138 => x"29810004",
    17139 => x"29630000", 17140 => x"b9a01000", 17141 => x"f8000199",
    17142 => x"5980000c", 17143 => x"59800008", 17144 => x"2b9d0004",
    17145 => x"2b8b0010", 17146 => x"2b8c000c", 17147 => x"2b8d0008",
    17148 => x"379c0010", 17149 => x"c3a00000", 17150 => x"379cfff8",
    17151 => x"5b8b0008", 17152 => x"5b9d0004", 17153 => x"b8205800",
    17154 => x"28210000", 17155 => x"f800016c", 17156 => x"78010001",
    17157 => x"38218f30", 17158 => x"28210000", 17159 => x"34020001",
    17160 => x"34030009", 17161 => x"58220004", 17162 => x"5963000c",
    17163 => x"78030001", 17164 => x"38635ab0", 17165 => x"59620008",
    17166 => x"28620000", 17167 => x"5822004c", 17168 => x"2b9d0004",
    17169 => x"2b8b0008", 17170 => x"379c0008", 17171 => x"c3a00000",
    17172 => x"b8201000", 17173 => x"28210000", 17174 => x"2823004c",
    17175 => x"34010000", 17176 => x"44600016", 17177 => x"28430004",
    17178 => x"28630038", 17179 => x"44600013", 17180 => x"78030001",
    17181 => x"38638f30", 17182 => x"28630000", 17183 => x"28640004",
    17184 => x"20840004", 17185 => x"4480000d", 17186 => x"28630004",
    17187 => x"20630008", 17188 => x"5c60000a", 17189 => x"2842000c",
    17190 => x"3403000a", 17191 => x"34010001", 17192 => x"54430006",
    17193 => x"78010001", 17194 => x"3c420002", 17195 => x"38215e8c",
    17196 => x"b4220800", 17197 => x"28210000", 17198 => x"c3a00000",
    17199 => x"379cfff0", 17200 => x"5b8b000c", 17201 => x"5b8c0008",
    17202 => x"5b9d0004", 17203 => x"2822000c", 17204 => x"b8205800",
    17205 => x"34010009", 17206 => x"3442ffff", 17207 => x"340c0000",
    17208 => x"544100a5", 17209 => x"78010001", 17210 => x"3c420002",
    17211 => x"38215e64", 17212 => x"b4220800", 17213 => x"28210000",
    17214 => x"c0200000", 17215 => x"78010001", 17216 => x"38218f30",
    17217 => x"28210000", 17218 => x"340c0000", 17219 => x"28220004",
    17220 => x"20420008", 17221 => x"5c400098", 17222 => x"28230004",
    17223 => x"78028000", 17224 => x"b8621000", 17225 => x"58220004",
    17226 => x"3401000a", 17227 => x"e0000090", 17228 => x"78010001",
    17229 => x"38218f30", 17230 => x"28210000", 17231 => x"78040001",
    17232 => x"38845a68", 17233 => x"28230004", 17234 => x"28820000",
    17235 => x"a0621000", 17236 => x"58220004", 17237 => x"28220004",
    17238 => x"20420008", 17239 => x"5c400083", 17240 => x"28210004",
    17241 => x"340c0001", 17242 => x"20210004", 17243 => x"44220082",
    17244 => x"596c000c", 17245 => x"e0000080", 17246 => x"29610000",
    17247 => x"340c0000", 17248 => x"2821004c", 17249 => x"4420007c",
    17250 => x"fbffbd10", 17251 => x"29610004", 17252 => x"f8000151",
    17253 => x"fbffbd16", 17254 => x"34010008", 17255 => x"e0000074",
    17256 => x"78010001", 17257 => x"38218f30", 17258 => x"28210000",
    17259 => x"34020002", 17260 => x"340c0000", 17261 => x"58220008",
    17262 => x"29610000", 17263 => x"2821004c", 17264 => x"4420006d",
    17265 => x"29610004", 17266 => x"28210038", 17267 => x"4420006a",
    17268 => x"78010001", 17269 => x"38218f44", 17270 => x"28210000",
    17271 => x"340300a2", 17272 => x"58230000", 17273 => x"34030003",
    17274 => x"58230010", 17275 => x"34030001", 17276 => x"5823001c",
    17277 => x"5962000c", 17278 => x"e000005e", 17279 => x"78010001",
    17280 => x"38218f44", 17281 => x"28210000", 17282 => x"340c0000",
    17283 => x"2822001c", 17284 => x"20420001", 17285 => x"44400058",
    17286 => x"34020002", 17287 => x"5822001c", 17288 => x"fbfff427",
    17289 => x"342107d0", 17290 => x"59610010", 17291 => x"34010003",
    17292 => x"e000004f", 17293 => x"fbfff422", 17294 => x"29620010",
    17295 => x"340c0000", 17296 => x"c8220800", 17297 => x"4801004c",
    17298 => x"34010007", 17299 => x"5961000c", 17300 => x"5960001c",
    17301 => x"e0000047", 17302 => x"37810010", 17303 => x"fbffff37",
    17304 => x"340c0000", 17305 => x"44200044", 17306 => x"78030001",
    17307 => x"38635ab4", 17308 => x"28620000", 17309 => x"2b810010",
    17310 => x"f80007a4", 17311 => x"3802c34f", 17312 => x"e8221000",
    17313 => x"64210000", 17314 => x"b8410800", 17315 => x"44200005",
    17316 => x"34010064", 17317 => x"59610014", 17318 => x"3401ff9c",
    17319 => x"e0000003", 17320 => x"59600014", 17321 => x"34010064",
    17322 => x"59610018", 17323 => x"34010004", 17324 => x"e000002f",
    17325 => x"29610004", 17326 => x"340c0000", 17327 => x"f80001df",
    17328 => x"5c20002d", 17329 => x"37810010", 17330 => x"fbffff1c",
    17331 => x"442c002a", 17332 => x"78040001", 17333 => x"38845ab4",
    17334 => x"2b810010", 17335 => x"28820000", 17336 => x"f800078a",
    17337 => x"29620014", 17338 => x"5b810010", 17339 => x"44220009",
    17340 => x"2961001c", 17341 => x"29620018", 17342 => x"b4410800",
    17343 => x"5961001c", 17344 => x"29610004", 17345 => x"2962001c",
    17346 => x"f80001aa", 17347 => x"e0000019", 17348 => x"29620014",
    17349 => x"340c0001", 17350 => x"5c220017", 17351 => x"2961001c",
    17352 => x"34217530", 17353 => x"5961001c", 17354 => x"29610004",
    17355 => x"2962001c", 17356 => x"f80001a0", 17357 => x"34010005",
    17358 => x"5961000c", 17359 => x"e000000e", 17360 => x"29610004",
    17361 => x"340c0000", 17362 => x"f80001bc", 17363 => x"5c20000a",
    17364 => x"34010006", 17365 => x"e0000006", 17366 => x"b9600800",
    17367 => x"fbffff3d", 17368 => x"340c0000", 17369 => x"5c200004",
    17370 => x"34010009", 17371 => x"5961000c", 17372 => x"340c0001",
    17373 => x"b9800800", 17374 => x"2b9d0004", 17375 => x"2b8b000c",
    17376 => x"2b8c0008", 17377 => x"379c0010", 17378 => x"c3a00000",
    17379 => x"78040001", 17380 => x"64630000", 17381 => x"38848f30",
    17382 => x"28850000", 17383 => x"c8031800", 17384 => x"78048000",
    17385 => x"78060001", 17386 => x"a0641800", 17387 => x"38c65ab8",
    17388 => x"b4641800", 17389 => x"28c40000", 17390 => x"3c210018",
    17391 => x"a0441000", 17392 => x"b8410800", 17393 => x"b8231800",
    17394 => x"58a3004c", 17395 => x"c3a00000", 17396 => x"78040001",
    17397 => x"64630000", 17398 => x"38848f30", 17399 => x"28850000",
    17400 => x"c8031800", 17401 => x"78048000", 17402 => x"78060001",
    17403 => x"a0641800", 17404 => x"38c65ab8", 17405 => x"b4641800",
    17406 => x"28c40000", 17407 => x"3c210018", 17408 => x"a0441000",
    17409 => x"b8410800", 17410 => x"b8231800", 17411 => x"58a3004c",
    17412 => x"c3a00000", 17413 => x"34030005", 17414 => x"5823002c",
    17415 => x"3803fffb", 17416 => x"58230030", 17417 => x"3403ff6a",
    17418 => x"5823001c", 17419 => x"3403fffe", 17420 => x"58230018",
    17421 => x"34030001", 17422 => x"58230028", 17423 => x"340300c8",
    17424 => x"58230048", 17425 => x"34032710", 17426 => x"58230040",
    17427 => x"34030064", 17428 => x"58230044", 17429 => x"5822000c",
    17430 => x"58200014", 17431 => x"c3a00000", 17432 => x"379cfff0",
    17433 => x"5b8b0010", 17434 => x"5b8c000c", 17435 => x"5b8d0008",
    17436 => x"5b9d0004", 17437 => x"b8205800", 17438 => x"2821000c",
    17439 => x"b8406800", 17440 => x"340c0000", 17441 => x"5c610047",
    17442 => x"34010022", 17443 => x"34030000", 17444 => x"fbffffbf",
    17445 => x"29620004", 17446 => x"34010025", 17447 => x"34030000",
    17448 => x"fbffffbb", 17449 => x"29610008", 17450 => x"4c200004",
    17451 => x"596d0004", 17452 => x"596d0008", 17453 => x"e000003b",
    17454 => x"4da10005", 17455 => x"29620000", 17456 => x"78010040",
    17457 => x"b4410800", 17458 => x"59610000", 17459 => x"29630000",
    17460 => x"78050001", 17461 => x"29620004", 17462 => x"38a55abc",
    17463 => x"28a10000", 17464 => x"b5a32000", 17465 => x"c8826000",
    17466 => x"482c0006", 17467 => x"78050001", 17468 => x"38a55ac0",
    17469 => x"28a10000", 17470 => x"49810002", 17471 => x"e0000002",
    17472 => x"b8206000", 17473 => x"78050001", 17474 => x"38a55ac4",
    17475 => x"28a10000", 17476 => x"4c240006", 17477 => x"4c220005",
    17478 => x"c8611800", 17479 => x"c8410800", 17480 => x"59630000",
    17481 => x"59610004", 17482 => x"29610004", 17483 => x"b9801000",
    17484 => x"596d0008", 17485 => x"34214000", 17486 => x"59610004",
    17487 => x"35610018", 17488 => x"fbfffdec", 17489 => x"78030001",
    17490 => x"38638f30", 17491 => x"29620010", 17492 => x"b8206800",
    17493 => x"28610000", 17494 => x"34030000", 17495 => x"582d0040",
    17496 => x"34410001", 17497 => x"59610010", 17498 => x"34010026",
    17499 => x"fbffff88", 17500 => x"34010020", 17501 => x"b9a01000",
    17502 => x"34030000", 17503 => x"fbffff84", 17504 => x"b9801000",
    17505 => x"34010021", 17506 => x"34030001", 17507 => x"fbffff80",
    17508 => x"b9801000", 17509 => x"3561003c", 17510 => x"fbfffdf7",
    17511 => x"7c2c0000", 17512 => x"b9800800", 17513 => x"2b9d0004",
    17514 => x"2b8b0010", 17515 => x"2b8c000c", 17516 => x"2b8d0008",
    17517 => x"379c0010", 17518 => x"c3a00000", 17519 => x"379cfff8",
    17520 => x"5b8b0008", 17521 => x"5b9d0004", 17522 => x"b8205800",
    17523 => x"2821002c", 17524 => x"59600004", 17525 => x"59600000",
    17526 => x"59610024", 17527 => x"3401ffff", 17528 => x"59610008",
    17529 => x"59600010", 17530 => x"35610018", 17531 => x"fbfffdde",
    17532 => x"3561003c", 17533 => x"fbfffe05", 17534 => x"78020001",
    17535 => x"35610054", 17536 => x"34030010", 17537 => x"38425eb8",
    17538 => x"fbfffe2b", 17539 => x"2961000c", 17540 => x"34020001",
    17541 => x"fbfffe01", 17542 => x"34010024", 17543 => x"34020001",
    17544 => x"34030001", 17545 => x"fbffff5a", 17546 => x"2b9d0004",
    17547 => x"2b8b0008", 17548 => x"379c0008", 17549 => x"c3a00000",
    17550 => x"379cfff8", 17551 => x"5b8b0008", 17552 => x"5b9d0004",
    17553 => x"b8205800", 17554 => x"34010005", 17555 => x"59610018",
    17556 => x"3801fffa", 17557 => x"5961001c", 17558 => x"34010001",
    17559 => x"59610014", 17560 => x"34017530", 17561 => x"59610010",
    17562 => x"3401fbb4", 17563 => x"59610008", 17564 => x"3401ffe2",
    17565 => x"59610004", 17566 => x"340104b0", 17567 => x"59610034",
    17568 => x"340103e8", 17569 => x"5961002c", 17570 => x"34010064",
    17571 => x"59610030", 17572 => x"78010001", 17573 => x"38219294",
    17574 => x"28210000", 17575 => x"59630074", 17576 => x"59620070",
    17577 => x"c8611800", 17578 => x"59630080", 17579 => x"35610004",
    17580 => x"5960007c", 17581 => x"59600084", 17582 => x"fbfffdab",
    17583 => x"35610028", 17584 => x"fbfffdd2", 17585 => x"2b9d0004",
    17586 => x"2b8b0008", 17587 => x"379c0008", 17588 => x"c3a00000",
    17589 => x"379cfff8", 17590 => x"5b8b0008", 17591 => x"5b9d0004",
    17592 => x"b8205800", 17593 => x"58200044", 17594 => x"58200040",
    17595 => x"3401ffff", 17596 => x"59610048", 17597 => x"5961004c",
    17598 => x"59610050", 17599 => x"59610054", 17600 => x"34010001",
    17601 => x"59610084", 17602 => x"59600058", 17603 => x"35610004",
    17604 => x"5960005c", 17605 => x"59600060", 17606 => x"59600068",
    17607 => x"5960006c", 17608 => x"59600078", 17609 => x"fbfffd90",
    17610 => x"35610028", 17611 => x"fbfffdb7", 17612 => x"29610070",
    17613 => x"34020001", 17614 => x"fbfffdb8", 17615 => x"29610074",
    17616 => x"34020001", 17617 => x"fbfffdb5", 17618 => x"34010004",
    17619 => x"34020001", 17620 => x"34030001", 17621 => x"fbffff1f",
    17622 => x"2b9d0004", 17623 => x"2b8b0008", 17624 => x"379c0008",
    17625 => x"c3a00000", 17626 => x"379cfff8", 17627 => x"5b8b0008",
    17628 => x"5b9d0004", 17629 => x"b8205800", 17630 => x"28210074",
    17631 => x"34020000", 17632 => x"fbfffda6", 17633 => x"59600084",
    17634 => x"2b9d0004", 17635 => x"2b8b0008", 17636 => x"379c0008",
    17637 => x"c3a00000", 17638 => x"379cfff0", 17639 => x"5b8b0010",
    17640 => x"5b8c000c", 17641 => x"5b8d0008", 17642 => x"5b9d0004",
    17643 => x"28240084", 17644 => x"b8205800", 17645 => x"34010001",
    17646 => x"44800078", 17647 => x"29610070", 17648 => x"5c610002",
    17649 => x"59620048", 17650 => x"29610074", 17651 => x"5c610002",
    17652 => x"5962004c", 17653 => x"29610048", 17654 => x"48010009",
    17655 => x"29620050", 17656 => x"48020006", 17657 => x"4c220005",
    17658 => x"29630040", 17659 => x"78020040", 17660 => x"b4621000",
    17661 => x"59620040", 17662 => x"59610050", 17663 => x"2961004c",
    17664 => x"48010009", 17665 => x"29620054", 17666 => x"48020006",
    17667 => x"4c220005", 17668 => x"29630044", 17669 => x"78020040",
    17670 => x"b4621000", 17671 => x"59620044", 17672 => x"59610054",
    17673 => x"29630048", 17674 => x"34010000", 17675 => x"4803005b",
    17676 => x"2962004c", 17677 => x"48020059", 17678 => x"296c0040",
    17679 => x"29610038", 17680 => x"b46c1800", 17681 => x"296c0044",
    17682 => x"c8621000", 17683 => x"c84c6000", 17684 => x"44200006",
    17685 => x"218c3fff", 17686 => x"21812000", 17687 => x"44200003",
    17688 => x"3401c000", 17689 => x"b9816000", 17690 => x"b9801000",
    17691 => x"35610004", 17692 => x"fbfffd20", 17693 => x"29620080",
    17694 => x"78030001", 17695 => x"38638f30", 17696 => x"2042000f",
    17697 => x"b8206800", 17698 => x"3c420010", 17699 => x"28610000",
    17700 => x"21a3ffff", 17701 => x"b8621000", 17702 => x"58220044",
    17703 => x"29630040", 17704 => x"29620048", 17705 => x"34010005",
    17706 => x"b4621000", 17707 => x"34030000", 17708 => x"fbfffec8",
    17709 => x"29630044", 17710 => x"2962004c", 17711 => x"34010002",
    17712 => x"b4621000", 17713 => x"34030000", 17714 => x"fbfffec2",
    17715 => x"34010001", 17716 => x"b9801000", 17717 => x"34030000",
    17718 => x"fbfffebe", 17719 => x"29620078", 17720 => x"34030000",
    17721 => x"34410001", 17722 => x"59610078", 17723 => x"34010006",
    17724 => x"fbfffeb8", 17725 => x"34010000", 17726 => x"b9a01000",
    17727 => x"34030001", 17728 => x"fbfffeb4", 17729 => x"78020001",
    17730 => x"3401ffff", 17731 => x"38425ac8", 17732 => x"5961004c",
    17733 => x"59610048", 17734 => x"29630040", 17735 => x"28410000",
    17736 => x"4c23000a", 17737 => x"29620044", 17738 => x"4c220008",
    17739 => x"78040001", 17740 => x"38845acc", 17741 => x"28810000",
    17742 => x"b4611800", 17743 => x"b4410800", 17744 => x"59630040",
    17745 => x"59610044", 17746 => x"29610038", 17747 => x"4420000f",
    17748 => x"2961006c", 17749 => x"29620068", 17750 => x"4c220006",
    17751 => x"34210001", 17752 => x"5961006c", 17753 => x"29610040",
    17754 => x"3421ffff", 17755 => x"e0000006", 17756 => x"4c410006",
    17757 => x"3421ffff", 17758 => x"5961006c", 17759 => x"29610040",
    17760 => x"34210001", 17761 => x"59610040", 17762 => x"35610028",
    17763 => x"b9801000", 17764 => x"fbfffcf9", 17765 => x"7c210000",
    17766 => x"2b9d0004", 17767 => x"2b8b0010", 17768 => x"2b8c000c",
    17769 => x"2b8d0008", 17770 => x"379c0010", 17771 => x"c3a00000",
    17772 => x"379cfff0", 17773 => x"5b8b0008", 17774 => x"5b9d0004",
    17775 => x"b8205800", 17776 => x"1443001f", 17777 => x"3781000c",
    17778 => x"4802000b", 17779 => x"00440012", 17780 => x"3c63000e",
    17781 => x"3c42000e", 17782 => x"b8641800", 17783 => x"5b820010",
    17784 => x"34021f40", 17785 => x"5b83000c", 17786 => x"fbffc100",
    17787 => x"2b820010", 17788 => x"e0000009", 17789 => x"0842c000",
    17790 => x"5b820010", 17791 => x"1442001f", 17792 => x"5b82000c",
    17793 => x"34021f40", 17794 => x"fbffc0f8", 17795 => x"2b820010",
    17796 => x"c8021000", 17797 => x"0041001f", 17798 => x"b4221000",
    17799 => x"14420001", 17800 => x"34010000", 17801 => x"59620068",
    17802 => x"2b9d0004", 17803 => x"2b8b0008", 17804 => x"379c0010",
    17805 => x"c3a00000", 17806 => x"28220068", 17807 => x"2821006c",
    17808 => x"fc410800", 17809 => x"c3a00000", 17810 => x"58220004",
    17811 => x"5820001c", 17812 => x"58230008", 17813 => x"5820000c",
    17814 => x"58200010", 17815 => x"58200000", 17816 => x"c3a00000",
    17817 => x"379cfffc", 17818 => x"5b9d0004", 17819 => x"34020001",
    17820 => x"58220000", 17821 => x"58200014", 17822 => x"5820001c",
    17823 => x"5820000c", 17824 => x"58200010", 17825 => x"28210004",
    17826 => x"fbfffce4", 17827 => x"78010001", 17828 => x"38219294",
    17829 => x"28210000", 17830 => x"34020001", 17831 => x"fbfffcdf",
    17832 => x"2b9d0004", 17833 => x"379c0004", 17834 => x"c3a00000",
    17835 => x"379cffb0", 17836 => x"5b8b0010", 17837 => x"5b8c000c",
    17838 => x"5b8d0008", 17839 => x"5b9d0004", 17840 => x"b8205800",
    17841 => x"b8406000", 17842 => x"b8606800", 17843 => x"37810014",
    17844 => x"34020000", 17845 => x"34030040", 17846 => x"f800068b",
    17847 => x"3401c000", 17848 => x"78040001", 17849 => x"5b810020",
    17850 => x"38849294", 17851 => x"34014000", 17852 => x"5b810044",
    17853 => x"28810000", 17854 => x"5da10005", 17855 => x"78030001",
    17856 => x"386372b4", 17857 => x"586c0000", 17858 => x"e0000027",
    17859 => x"3dad0005", 17860 => x"b56d5800", 17861 => x"29610000",
    17862 => x"44200023", 17863 => x"78030001", 17864 => x"386372b4",
    17865 => x"28610000", 17866 => x"29620010", 17867 => x"c9810800",
    17868 => x"20213fff", 17869 => x"1423000c", 17870 => x"5c400007",
    17871 => x"3c630002", 17872 => x"5961000c", 17873 => x"34010001",
    17874 => x"59630014", 17875 => x"59610010", 17876 => x"e0000015",
    17877 => x"2964000c", 17878 => x"34420001", 17879 => x"b4240800",
    17880 => x"29640014", 17881 => x"b4641800", 17882 => x"3c630002",
    17883 => x"37840050", 17884 => x"b4831800", 17885 => x"2863ffc4",
    17886 => x"59620010", 17887 => x"b4230800", 17888 => x"29630008",
    17889 => x"5961000c", 17890 => x"5c430007", 17891 => x"f8000532",
    17892 => x"59610018", 17893 => x"34010001", 17894 => x"5961001c",
    17895 => x"5960000c", 17896 => x"59600010", 17897 => x"34010000",
    17898 => x"2b9d0004", 17899 => x"2b8b0010", 17900 => x"2b8c000c",
    17901 => x"2b8d0008", 17902 => x"379c0050", 17903 => x"c3a00000",
    17904 => x"78030001", 17905 => x"38638f30", 17906 => x"5c40000a",
    17907 => x"34040001", 17908 => x"28620000", 17909 => x"bc810800",
    17910 => x"202100ff", 17911 => x"28430020", 17912 => x"3c210010",
    17913 => x"a4200800", 17914 => x"a0230800", 17915 => x"e0000008",
    17916 => x"28620000", 17917 => x"34040001", 17918 => x"bc810800",
    17919 => x"28430020", 17920 => x"202100ff", 17921 => x"3c210010",
    17922 => x"b8230800", 17923 => x"58410020", 17924 => x"c3a00000",
    17925 => x"379cfff8", 17926 => x"5b8b0008", 17927 => x"5b9d0004",
    17928 => x"34020001", 17929 => x"44220009", 17930 => x"34020002",
    17931 => x"4422000c", 17932 => x"5c200017", 17933 => x"78010001",
    17934 => x"38218f30", 17935 => x"282b0000", 17936 => x"356b0018",
    17937 => x"e000000a", 17938 => x"78010001", 17939 => x"38218f30",
    17940 => x"282b0000", 17941 => x"356b0014", 17942 => x"e0000005",
    17943 => x"78010001", 17944 => x"38218f30", 17945 => x"282b0000",
    17946 => x"356b001c", 17947 => x"340107d0", 17948 => x"fbfff198",
    17949 => x"78030001", 17950 => x"38635a88", 17951 => x"29620000",
    17952 => x"28610000", 17953 => x"a0410800", 17954 => x"e0000002",
    17955 => x"34010000", 17956 => x"2b9d0004", 17957 => x"2b8b0008",
    17958 => x"379c0008", 17959 => x"c3a00000", 17960 => x"379cfff8",
    17961 => x"5b8b0008", 17962 => x"5b9d0004", 17963 => x"b8201800",
    17964 => x"78010001", 17965 => x"b8405800", 17966 => x"38219004",
    17967 => x"44600007", 17968 => x"3461ffff", 17969 => x"08210090",
    17970 => x"78030001", 17971 => x"38638f4c", 17972 => x"34210148",
    17973 => x"b4230800", 17974 => x"b9601000", 17975 => x"fbffff35",
    17976 => x"78010001", 17977 => x"38218f4c", 17978 => x"582b0018",
    17979 => x"2b9d0004", 17980 => x"2b8b0008", 17981 => x"379c0008",
    17982 => x"c3a00000", 17983 => x"379cffec", 17984 => x"5b8b0014",
    17985 => x"5b8c0010", 17986 => x"5b8d000c", 17987 => x"5b8e0008",
    17988 => x"5b9d0004", 17989 => x"780c0001", 17990 => x"780d0001",
    17991 => x"b8207000", 17992 => x"340b0000", 17993 => x"398c9294",
    17994 => x"39ad8f20", 17995 => x"e000000a", 17996 => x"29a10000",
    17997 => x"942b0800", 17998 => x"20210001", 17999 => x"44200005",
    18000 => x"35620013", 18001 => x"3c420005", 18002 => x"b5c20800",
    18003 => x"fbffff46", 18004 => x"356b0001", 18005 => x"29810000",
    18006 => x"482bfff6", 18007 => x"2b9d0004", 18008 => x"2b8b0014",
    18009 => x"2b8c0010", 18010 => x"2b8d000c", 18011 => x"2b8e0008",
    18012 => x"379c0014", 18013 => x"c3a00000", 18014 => x"379cffbc",
    18015 => x"5b8b0044", 18016 => x"5b8c0040", 18017 => x"5b8d003c",
    18018 => x"5b8e0038", 18019 => x"5b8f0034", 18020 => x"5b900030",
    18021 => x"5b91002c", 18022 => x"5b920028", 18023 => x"5b930024",
    18024 => x"5b940020", 18025 => x"5b95001c", 18026 => x"5b960018",
    18027 => x"5b970014", 18028 => x"5b980010", 18029 => x"5b99000c",
    18030 => x"5b9b0008", 18031 => x"5b9d0004", 18032 => x"781b0001",
    18033 => x"780b0001", 18034 => x"78190001", 18035 => x"780d0001",
    18036 => x"78110001", 18037 => x"78100001", 18038 => x"780c0001",
    18039 => x"78170001", 18040 => x"780f0001", 18041 => x"3b7b8f30",
    18042 => x"396b8f4c", 18043 => x"34140009", 18044 => x"3b395ecc",
    18045 => x"34180001", 18046 => x"34130003", 18047 => x"39ad8fe4",
    18048 => x"34120008", 18049 => x"3a319004", 18050 => x"3a108f68",
    18051 => x"398c9294", 18052 => x"3af791ac", 18053 => x"39ef928c",
    18054 => x"e0000079", 18055 => x"2875007c", 18056 => x"780100ff",
    18057 => x"3821ffff", 18058 => x"02ae0018", 18059 => x"a2a1a800",
    18060 => x"29610004", 18061 => x"21ce007f", 18062 => x"3421ffff",
    18063 => x"54340050", 18064 => x"3c210002", 18065 => x"b7210800",
    18066 => x"28210000", 18067 => x"c0200000", 18068 => x"2961004c",
    18069 => x"58610040", 18070 => x"296100d4", 18071 => x"296200d0",
    18072 => x"b4410800", 18073 => x"0022001f", 18074 => x"b4410800",
    18075 => x"14210001", 18076 => x"34020001", 18077 => x"58610044",
    18078 => x"29810000", 18079 => x"fbfffbe7", 18080 => x"fbfff10f",
    18081 => x"34210032", 18082 => x"59610008", 18083 => x"3401000a",
    18084 => x"e0000011", 18085 => x"29760008", 18086 => x"fbfff109",
    18087 => x"cac10800", 18088 => x"4c200037", 18089 => x"29610000",
    18090 => x"5c380003", 18091 => x"59780004", 18092 => x"e0000033",
    18093 => x"59730004", 18094 => x"e0000031", 18095 => x"29810000",
    18096 => x"34020000", 18097 => x"fbfffbd5", 18098 => x"b9a00800",
    18099 => x"fbfffc4b", 18100 => x"34010002", 18101 => x"59610004",
    18102 => x"e0000029", 18103 => x"b9a00800", 18104 => x"fbfffc5c",
    18105 => x"e0000012", 18106 => x"ba000800", 18107 => x"fbfffdb4",
    18108 => x"34010004", 18109 => x"e3fffff8", 18110 => x"29610068",
    18111 => x"44200020", 18112 => x"2961006c", 18113 => x"4420001e",
    18114 => x"29610000", 18115 => x"5c330009", 18116 => x"34010005",
    18117 => x"e3fffff0", 18118 => x"ba200800", 18119 => x"fbfffdee",
    18120 => x"34010006", 18121 => x"e3ffffec", 18122 => x"296100f0",
    18123 => x"44200014", 18124 => x"b9600800", 18125 => x"fbffff72",
    18126 => x"59720004", 18127 => x"e0000010", 18128 => x"29610000",
    18129 => x"5c380004", 18130 => x"b9a00800", 18131 => x"fbfffc41",
    18132 => x"44200007", 18133 => x"29610068", 18134 => x"44200005",
    18135 => x"29610000", 18136 => x"5c330007", 18137 => x"296100f0",
    18138 => x"5c200005", 18139 => x"29610010", 18140 => x"34210001",
    18141 => x"59610010", 18142 => x"59740004", 18143 => x"ba000800",
    18144 => x"baa01000", 18145 => x"b9c01800", 18146 => x"fbfffd36",
    18147 => x"29610068", 18148 => x"4420001b", 18149 => x"ba200800",
    18150 => x"baa01000", 18151 => x"b9c01800", 18152 => x"fbfffdfe",
    18153 => x"29610004", 18154 => x"5c320015", 18155 => x"29610000",
    18156 => x"34160000", 18157 => x"5c33000c", 18158 => x"e0000008",
    18159 => x"0ac10090", 18160 => x"baa01000", 18161 => x"b9c01800",
    18162 => x"34210148", 18163 => x"b5610800", 18164 => x"fbfffdf2",
    18165 => x"36d60001", 18166 => x"29e10000", 18167 => x"3421ffff",
    18168 => x"4836fff7", 18169 => x"29810000", 18170 => x"49c10005",
    18171 => x"bae00800", 18172 => x"baa01000", 18173 => x"b9c01800",
    18174 => x"fbfffead", 18175 => x"2b630000", 18176 => x"78020002",
    18177 => x"28610080", 18178 => x"a0220800", 18179 => x"4420ff84",
    18180 => x"29610014", 18181 => x"34210001", 18182 => x"59610014",
    18183 => x"34010001", 18184 => x"d0410000", 18185 => x"2b9d0004",
    18186 => x"2b8b0044", 18187 => x"2b8c0040", 18188 => x"2b8d003c",
    18189 => x"2b8e0038", 18190 => x"2b8f0034", 18191 => x"2b900030",
    18192 => x"2b91002c", 18193 => x"2b920028", 18194 => x"2b930024",
    18195 => x"2b940020", 18196 => x"2b95001c", 18197 => x"2b960018",
    18198 => x"2b970014", 18199 => x"2b980010", 18200 => x"2b99000c",
    18201 => x"2b9b0008", 18202 => x"379c0044", 18203 => x"c3a00000",
    18204 => x"78010001", 18205 => x"38218f48", 18206 => x"28220000",
    18207 => x"78030001", 18208 => x"78010001", 18209 => x"38218f44",
    18210 => x"38635ad0", 18211 => x"58220000", 18212 => x"28610000",
    18213 => x"58410000", 18214 => x"c3a00000", 18215 => x"379cffd4",
    18216 => x"5b8b0028", 18217 => x"5b8c0024", 18218 => x"5b8d0020",
    18219 => x"5b8e001c", 18220 => x"5b8f0018", 18221 => x"5b900014",
    18222 => x"5b910010", 18223 => x"5b92000c", 18224 => x"5b930008",
    18225 => x"5b9d0004", 18226 => x"b8205800", 18227 => x"b8408000",
    18228 => x"b8609000", 18229 => x"fbffb93d", 18230 => x"78010001",
    18231 => x"382192c4", 18232 => x"28240000", 18233 => x"78010001",
    18234 => x"38218f30", 18235 => x"58240000", 18236 => x"78010001",
    18237 => x"28850000", 18238 => x"38218f48", 18239 => x"28210000",
    18240 => x"78020001", 18241 => x"38428f44", 18242 => x"00a60010",
    18243 => x"58410000", 18244 => x"78020001", 18245 => x"38429294",
    18246 => x"20c6003f", 18247 => x"00a50018", 18248 => x"58460000",
    18249 => x"78020001", 18250 => x"3842928c", 18251 => x"20a50007",
    18252 => x"58450000", 18253 => x"78050001", 18254 => x"38a58f4c",
    18255 => x"58ab0000", 18256 => x"58a00010", 18257 => x"58800040",
    18258 => x"58800044", 18259 => x"58800000", 18260 => x"58800028",
    18261 => x"58800024", 18262 => x"58800004", 18263 => x"78030001",
    18264 => x"58800020", 18265 => x"340203e8", 18266 => x"38635a9c",
    18267 => x"58820048", 18268 => x"28620000", 18269 => x"5820001c",
    18270 => x"58220000", 18271 => x"34010004", 18272 => x"5d610004",
    18273 => x"34010007", 18274 => x"58a10004", 18275 => x"e0000006",
    18276 => x"34010009", 18277 => x"58a10004", 18278 => x"34010003",
    18279 => x"5d610002", 18280 => x"ba003000", 18281 => x"78010001",
    18282 => x"b8c01000", 18283 => x"38218f68", 18284 => x"780d0001",
    18285 => x"fbfffc98", 18286 => x"39ad9294", 18287 => x"29a30000",
    18288 => x"78010001", 18289 => x"38219004", 18290 => x"ba001000",
    18291 => x"780f0001", 18292 => x"780e0001", 18293 => x"fbfffd19",
    18294 => x"340c0000", 18295 => x"39ef928c", 18296 => x"39ce8f4c",
    18297 => x"34130001", 18298 => x"e000000c", 18299 => x"09910090",
    18300 => x"29a40000", 18301 => x"ba001000", 18302 => x"36210148",
    18303 => x"34840001", 18304 => x"b48c1800", 18305 => x"b5c10800",
    18306 => x"b5d18800", 18307 => x"fbfffd0b", 18308 => x"358c0001",
    18309 => x"5a330140", 18310 => x"29e10000", 18311 => x"3421ffff",
    18312 => x"482cfff3", 18313 => x"34010002", 18314 => x"5d610006",
    18315 => x"78010001", 18316 => x"38218f44", 18317 => x"28210000",
    18318 => x"34020006", 18319 => x"5822001c", 18320 => x"780e0001",
    18321 => x"780d0001", 18322 => x"340c0000", 18323 => x"39ce9294",
    18324 => x"39ad8f4c", 18325 => x"e0000008", 18326 => x"35810013",
    18327 => x"3c210005", 18328 => x"b9801000", 18329 => x"b5a10800",
    18330 => x"34030200", 18331 => x"fbfffdf7", 18332 => x"358c0001",
    18333 => x"29c20000", 18334 => x"484cfff8", 18335 => x"34010001",
    18336 => x"5d610017", 18337 => x"78010001", 18338 => x"38218f30",
    18339 => x"28210000", 18340 => x"28210004", 18341 => x"20210002",
    18342 => x"44200021", 18343 => x"78010001", 18344 => x"78040001",
    18345 => x"38218f4c", 18346 => x"38848f68", 18347 => x"58240098",
    18348 => x"78040001", 18349 => x"38849004", 18350 => x"5824009c",
    18351 => x"78010001", 18352 => x"3821928c", 18353 => x"28240000",
    18354 => x"78010001", 18355 => x"38218fe4", 18356 => x"b4441000",
    18357 => x"ba401800", 18358 => x"fbfffb2c", 18359 => x"78010001",
    18360 => x"38218f30", 18361 => x"28210000", 18362 => x"78020002",
    18363 => x"e0000003", 18364 => x"2823007c", 18365 => x"5b83002c",
    18366 => x"28230080", 18367 => x"a0621800", 18368 => x"4460fffc",
    18369 => x"34020001", 18370 => x"58220064", 18371 => x"28220028",
    18372 => x"38420001", 18373 => x"58220028", 18374 => x"fbffb8b5",
    18375 => x"2b9d0004", 18376 => x"2b8b0028", 18377 => x"2b8c0024",
    18378 => x"2b8d0020", 18379 => x"2b8e001c", 18380 => x"2b8f0018",
    18381 => x"2b900014", 18382 => x"2b910010", 18383 => x"2b92000c",
    18384 => x"2b930008", 18385 => x"379c002c", 18386 => x"c3a00000",
    18387 => x"379cfffc", 18388 => x"5b9d0004", 18389 => x"78020001",
    18390 => x"38428f4c", 18391 => x"28430004", 18392 => x"64240000",
    18393 => x"7c630008", 18394 => x"b8831800", 18395 => x"5c600006",
    18396 => x"3421ffff", 18397 => x"08210090", 18398 => x"34210148",
    18399 => x"b4410800", 18400 => x"fbfffcd5", 18401 => x"2b9d0004",
    18402 => x"379c0004", 18403 => x"c3a00000", 18404 => x"379cfffc",
    18405 => x"5b9d0004", 18406 => x"44200008", 18407 => x"3421ffff",
    18408 => x"08210090", 18409 => x"78020001", 18410 => x"38428f4c",
    18411 => x"34210148", 18412 => x"b4220800", 18413 => x"fbfffced",
    18414 => x"2b9d0004", 18415 => x"379c0004", 18416 => x"c3a00000",
    18417 => x"78020001", 18418 => x"b8201800", 18419 => x"38428f4c",
    18420 => x"5c200004", 18421 => x"28410004", 18422 => x"64210008",
    18423 => x"c3a00000", 18424 => x"28450004", 18425 => x"34040008",
    18426 => x"34010000", 18427 => x"5ca40006", 18428 => x"3463ffff",
    18429 => x"08630090", 18430 => x"b4431000", 18431 => x"28410180",
    18432 => x"7c210000", 18433 => x"c3a00000", 18434 => x"379cffe8",
    18435 => x"5b8b0018", 18436 => x"5b8c0014", 18437 => x"5b8d0010",
    18438 => x"5b8e000c", 18439 => x"5b8f0008", 18440 => x"5b9d0004",
    18441 => x"3403ffff", 18442 => x"b8407800", 18443 => x"5c230016",
    18444 => x"34010000", 18445 => x"780c0001", 18446 => x"780d0001",
    18447 => x"fbfffe19", 18448 => x"340b0000", 18449 => x"398c928c",
    18450 => x"39ad8f4c", 18451 => x"340e0004", 18452 => x"e0000009",
    18453 => x"09610090", 18454 => x"b5a10800", 18455 => x"28210140",
    18456 => x"5c2e0004", 18457 => x"35610001", 18458 => x"b9e01000",
    18459 => x"fbfffe0d", 18460 => x"356b0001", 18461 => x"29810000",
    18462 => x"3421ffff", 18463 => x"482bfff6", 18464 => x"e0000002",
    18465 => x"fbfffe07", 18466 => x"2b9d0004", 18467 => x"2b8b0018",
    18468 => x"2b8c0014", 18469 => x"2b8d0010", 18470 => x"2b8e000c",
    18471 => x"2b8f0008", 18472 => x"379c0018", 18473 => x"c3a00000",
    18474 => x"379cfff0", 18475 => x"5b8b0010", 18476 => x"5b8c000c",
    18477 => x"5b8d0008", 18478 => x"5b9d0004", 18479 => x"780b0001",
    18480 => x"b8406800", 18481 => x"b8606000", 18482 => x"396b9004",
    18483 => x"44200007", 18484 => x"342bffff", 18485 => x"096b0090",
    18486 => x"78010001", 18487 => x"38218f4c", 18488 => x"356b0148",
    18489 => x"b5615800", 18490 => x"45a0000b", 18491 => x"2962006c",
    18492 => x"34041f40", 18493 => x"34030000", 18494 => x"3c420001",
    18495 => x"1441001f", 18496 => x"f80002ae", 18497 => x"3c210012",
    18498 => x"0044000e", 18499 => x"b8242000", 18500 => x"59a40000",
    18501 => x"4580000b", 18502 => x"29620068", 18503 => x"34030000",
    18504 => x"34041f40", 18505 => x"3c420001", 18506 => x"1441001f",
    18507 => x"f80002a3", 18508 => x"3c210012", 18509 => x"0042000e",
    18510 => x"b8221000", 18511 => x"59820000", 18512 => x"2b9d0004",
    18513 => x"2b8b0010", 18514 => x"2b8c000c", 18515 => x"2b8d0008",
    18516 => x"379c0010", 18517 => x"c3a00000", 18518 => x"379cfff0",
    18519 => x"5b8b0010", 18520 => x"5b8c000c", 18521 => x"5b8d0008",
    18522 => x"5b9d0004", 18523 => x"b8205800", 18524 => x"b8406800",
    18525 => x"78010001", 18526 => x"3d620005", 18527 => x"38218f4c",
    18528 => x"b4220800", 18529 => x"28240278", 18530 => x"b8606000",
    18531 => x"4c800003", 18532 => x"34844000", 18533 => x"e0000004",
    18534 => x"34013fff", 18535 => x"4c240002", 18536 => x"3484c000",
    18537 => x"3c840001", 18538 => x"34010000", 18539 => x"20823ffe",
    18540 => x"34030000", 18541 => x"34041f40", 18542 => x"f8000280",
    18543 => x"3c210012", 18544 => x"0044000e", 18545 => x"b8242000",
    18546 => x"59a40000", 18547 => x"4580000d", 18548 => x"78010001",
    18549 => x"38218f20", 18550 => x"35630013", 18551 => x"28220000",
    18552 => x"3c630005", 18553 => x"78010001", 18554 => x"38218f4c",
    18555 => x"b4230800", 18556 => x"28210004", 18557 => x"94410800",
    18558 => x"20210001", 18559 => x"59810000", 18560 => x"3d6b0005",
    18561 => x"78020001", 18562 => x"38428f4c", 18563 => x"b44b1000",
    18564 => x"2841027c", 18565 => x"2b9d0004", 18566 => x"2b8b0010",
    18567 => x"2b8c000c", 18568 => x"2b8d0008", 18569 => x"379c0010",
    18570 => x"c3a00000", 18571 => x"379cffec", 18572 => x"5b8b0014",
    18573 => x"5b8c0010", 18574 => x"5b9d000c", 18575 => x"780b0001",
    18576 => x"396b8f4c", 18577 => x"29610000", 18578 => x"4c010014",
    18579 => x"296c0014", 18580 => x"29620004", 18581 => x"78010001",
    18582 => x"38215ef4", 18583 => x"fbfffa2c", 18584 => x"29640000",
    18585 => x"b8201800", 18586 => x"296500a4", 18587 => x"29660068",
    18588 => x"296700f0", 18589 => x"29680054", 18590 => x"296200dc",
    18591 => x"29610010", 18592 => x"5b820004", 18593 => x"5b810008",
    18594 => x"78010001", 18595 => x"38215950", 18596 => x"b9801000",
    18597 => x"fbffe94a", 18598 => x"2b9d000c", 18599 => x"2b8b0014",
    18600 => x"2b8c0010", 18601 => x"379c0014", 18602 => x"c3a00000",
    18603 => x"379cfffc", 18604 => x"5b9d0004", 18605 => x"5c200004",
    18606 => x"78010001", 18607 => x"38219004", 18608 => x"e0000007",
    18609 => x"3421ffff", 18610 => x"08210090", 18611 => x"78020001",
    18612 => x"38428f4c", 18613 => x"34210148", 18614 => x"b4220800",
    18615 => x"fbfffcd7", 18616 => x"2b9d0004", 18617 => x"379c0004",
    18618 => x"c3a00000", 18619 => x"379cfff0", 18620 => x"5b8b0010",
    18621 => x"5b8c000c", 18622 => x"5b8d0008", 18623 => x"5b9d0004",
    18624 => x"780d0001", 18625 => x"780b0001", 18626 => x"b8206000",
    18627 => x"39ad8f4c", 18628 => x"396b8f20", 18629 => x"4440000d",
    18630 => x"34020001", 18631 => x"fbfff9bf", 18632 => x"35810013",
    18633 => x"3c210005", 18634 => x"b5a10800", 18635 => x"fbfffcce",
    18636 => x"29610000", 18637 => x"34020001", 18638 => x"bc4c6000",
    18639 => x"b9816000", 18640 => x"596c0000", 18641 => x"e000000a",
    18642 => x"34030001", 18643 => x"29640000", 18644 => x"bc611800",
    18645 => x"a4601800", 18646 => x"a0641800", 18647 => x"59630000",
    18648 => x"29a30128", 18649 => x"44230002", 18650 => x"fbfff9ac",
    18651 => x"2b9d0004", 18652 => x"2b8b0010", 18653 => x"2b8c000c",
    18654 => x"2b8d0008", 18655 => x"379c0010", 18656 => x"c3a00000",
    18657 => x"08210090", 18658 => x"78020001", 18659 => x"38428f4c",
    18660 => x"b4411000", 18661 => x"28410140", 18662 => x"28430140",
    18663 => x"34020004", 18664 => x"7c210001", 18665 => x"5c620002",
    18666 => x"38210002", 18667 => x"c3a00000", 18668 => x"4c200005",
    18669 => x"78010001", 18670 => x"38218f4c", 18671 => x"28210054",
    18672 => x"c3a00000", 18673 => x"78020001", 18674 => x"38428f4c",
    18675 => x"5c200003", 18676 => x"284100dc", 18677 => x"c3a00000",
    18678 => x"3421ffff", 18679 => x"08210090", 18680 => x"b4411000",
    18681 => x"2841016c", 18682 => x"c3a00000", 18683 => x"78030001",
    18684 => x"38638f30", 18685 => x"4c200007", 18686 => x"78010001",
    18687 => x"38218f4c", 18688 => x"58220054", 18689 => x"28610000",
    18690 => x"58220040", 18691 => x"c3a00000", 18692 => x"2024000f",
    18693 => x"28630000", 18694 => x"3c840010", 18695 => x"2045ffff",
    18696 => x"b8a42000", 18697 => x"58640044", 18698 => x"78030001",
    18699 => x"38638f4c", 18700 => x"5c200003", 18701 => x"586200dc",
    18702 => x"c3a00000", 18703 => x"3421ffff", 18704 => x"08210090",
    18705 => x"b4611800", 18706 => x"5862016c", 18707 => x"c3a00000",
    18708 => x"379cffcc", 18709 => x"5b8b0034", 18710 => x"5b8c0030",
    18711 => x"5b8d002c", 18712 => x"5b8e0028", 18713 => x"5b8f0024",
    18714 => x"5b900020", 18715 => x"5b91001c", 18716 => x"5b920018",
    18717 => x"5b930014", 18718 => x"5b940010", 18719 => x"5b95000c",
    18720 => x"5b960008", 18721 => x"5b9d0004", 18722 => x"78010001",
    18723 => x"38218f4c", 18724 => x"28220000", 18725 => x"34010001",
    18726 => x"34140000", 18727 => x"5c410005", 18728 => x"78010001",
    18729 => x"38218fe4", 18730 => x"fbfffa05", 18731 => x"b820a000",
    18732 => x"78110001", 18733 => x"780b0001", 18734 => x"780e0001",
    18735 => x"340d0000", 18736 => x"340c0001", 18737 => x"3a31928c",
    18738 => x"396b8f4c", 18739 => x"340f0001", 18740 => x"39ce8f30",
    18741 => x"34120002", 18742 => x"34160003", 18743 => x"34150004",
    18744 => x"e0000047", 18745 => x"3593ffff", 18746 => x"0a700090",
    18747 => x"b5708000", 18748 => x"2a010140", 18749 => x"442f000f",
    18750 => x"29c10000", 18751 => x"bdec1000", 18752 => x"28210020",
    18753 => x"00210008", 18754 => x"202100ff", 18755 => x"a0220800",
    18756 => x"5c200008", 18757 => x"b9800800", 18758 => x"fbfffe9e",
    18759 => x"b9800800", 18760 => x"34020000", 18761 => x"fbfffca7",
    18762 => x"35ad0001", 18763 => x"5a0f0140", 18764 => x"0a610090",
    18765 => x"b5618000", 18766 => x"2a020140", 18767 => x"44520014",
    18768 => x"48520003", 18769 => x"5c4f002d", 18770 => x"e0000004",
    18771 => x"44560017", 18772 => x"5c55002a", 18773 => x"e000001e",
    18774 => x"296100f0", 18775 => x"44200027", 18776 => x"29c10000",
    18777 => x"bdec1000", 18778 => x"28210020", 18779 => x"00210008",
    18780 => x"202100ff", 18781 => x"a0220800", 18782 => x"44200020",
    18783 => x"b9800800", 18784 => x"fbfffe73", 18785 => x"5a120140",
    18786 => x"e000001b", 18787 => x"2a010180", 18788 => x"4420001a",
    18789 => x"29620018", 18790 => x"b9800800", 18791 => x"fbfffcc1",
    18792 => x"5a160140", 18793 => x"e0000014", 18794 => x"34210148",
    18795 => x"b5610800", 18796 => x"fbfffc22", 18797 => x"5c200011",
    18798 => x"b9800800", 18799 => x"34020001", 18800 => x"fbfffc80",
    18801 => x"5a150140", 18802 => x"e000000b", 18803 => x"296100f0",
    18804 => x"44200003", 18805 => x"2a010180", 18806 => x"5c200008",
    18807 => x"0a730090", 18808 => x"b9800800", 18809 => x"34020000",
    18810 => x"b5739800", 18811 => x"fbfffc75", 18812 => x"5a6f0140",
    18813 => x"35ad0001", 18814 => x"358c0001", 18815 => x"2a210000",
    18816 => x"482cffb9", 18817 => x"29630000", 18818 => x"78020001",
    18819 => x"384272bc", 18820 => x"5843000c", 18821 => x"29630014",
    18822 => x"28410008", 18823 => x"7dad0000", 18824 => x"58430010",
    18825 => x"29630004", 18826 => x"34210002", 18827 => x"b5b4a000",
    18828 => x"58430014", 18829 => x"296300a4", 18830 => x"58410008",
    18831 => x"7e810000", 18832 => x"58430018", 18833 => x"29630068",
    18834 => x"5843001c", 18835 => x"296300f0", 18836 => x"58430020",
    18837 => x"29630054", 18838 => x"58430024", 18839 => x"296300dc",
    18840 => x"58430028", 18841 => x"29630010", 18842 => x"5843002c",
    18843 => x"2b9d0004", 18844 => x"2b8b0034", 18845 => x"2b8c0030",
    18846 => x"2b8d002c", 18847 => x"2b8e0028", 18848 => x"2b8f0024",
    18849 => x"2b900020", 18850 => x"2b91001c", 18851 => x"2b920018",
    18852 => x"2b930014", 18853 => x"2b940010", 18854 => x"2b95000c",
    18855 => x"2b960008", 18856 => x"379c0034", 18857 => x"c3a00000",
    18858 => x"379cfff8", 18859 => x"5b8b0008", 18860 => x"5b9d0004",
    18861 => x"fbffb6c5", 18862 => x"34020000", 18863 => x"3401ffff",
    18864 => x"fbffff4b", 18865 => x"34010001", 18866 => x"fbfffc53",
    18867 => x"380bffff", 18868 => x"b9601000", 18869 => x"3401ffff",
    18870 => x"fbffff45", 18871 => x"34010001", 18872 => x"fbfffc4d",
    18873 => x"34020000", 18874 => x"34010000", 18875 => x"fbffff40",
    18876 => x"34010000", 18877 => x"fbfffc48", 18878 => x"b9601000",
    18879 => x"34010000", 18880 => x"fbffff3b", 18881 => x"34010000",
    18882 => x"fbfffc43", 18883 => x"34010002", 18884 => x"fbfffc41",
    18885 => x"2b9d0004", 18886 => x"2b8b0008", 18887 => x"379c0008",
    18888 => x"c3a00000", 18889 => x"379cfff0", 18890 => x"5b8b0010",
    18891 => x"5b8c000c", 18892 => x"5b8d0008", 18893 => x"5b9d0004",
    18894 => x"78010001", 18895 => x"780b0001", 18896 => x"38215a28",
    18897 => x"780c0001", 18898 => x"396bf800", 18899 => x"282d0000",
    18900 => x"398c5a14", 18901 => x"e0000005", 18902 => x"b9800800",
    18903 => x"fbffe818", 18904 => x"340103e8", 18905 => x"fbffeddb",
    18906 => x"29610000", 18907 => x"5c2dfffb", 18908 => x"2b9d0004",
    18909 => x"2b8b0010", 18910 => x"2b8c000c", 18911 => x"2b8d0008",
    18912 => x"379c0010", 18913 => x"c3a00000", 18914 => x"c3a00000",
    18915 => x"379cfff8", 18916 => x"5b8b0008", 18917 => x"5b9d0004",
    18918 => x"28240014", 18919 => x"b8201800", 18920 => x"b8403000",
    18921 => x"44800015", 18922 => x"28250010", 18923 => x"20a50002",
    18924 => x"5ca00007", 18925 => x"b4862000", 18926 => x"b8800800",
    18927 => x"2b9d0004", 18928 => x"2b8b0008", 18929 => x"379c0008",
    18930 => x"c3a00000", 18931 => x"346b0030", 18932 => x"b4861000",
    18933 => x"b9600800", 18934 => x"34030040", 18935 => x"f80001cc",
    18936 => x"b9602000", 18937 => x"b8800800", 18938 => x"2b9d0004",
    18939 => x"2b8b0008", 18940 => x"379c0008", 18941 => x"c3a00000",
    18942 => x"28250010", 18943 => x"20a70004", 18944 => x"5ce4ffeb",
    18945 => x"2825001c", 18946 => x"34040000", 18947 => x"44a7ffeb",
    18948 => x"342b0030", 18949 => x"34040040", 18950 => x"b9601800",
    18951 => x"d8a00000", 18952 => x"b9602000", 18953 => x"e3fffff0",
    18954 => x"379cfff4", 18955 => x"5b8b0008", 18956 => x"5b9d0004",
    18957 => x"28220014", 18958 => x"b8205800", 18959 => x"44400013",
    18960 => x"2961000c", 18961 => x"b4411000", 18962 => x"28430000",
    18963 => x"78040001", 18964 => x"38845ad4", 18965 => x"28820000",
    18966 => x"3401ffec", 18967 => x"5c620007", 18968 => x"78020001",
    18969 => x"38428f24", 18970 => x"28430000", 18971 => x"34010000",
    18972 => x"584b0000", 18973 => x"5963007c", 18974 => x"2b9d0004",
    18975 => x"2b8b0008", 18976 => x"379c000c", 18977 => x"c3a00000",
    18978 => x"28230010", 18979 => x"20630004", 18980 => x"5c62ffec",
    18981 => x"2825001c", 18982 => x"2822000c", 18983 => x"3783000c",
    18984 => x"34040004", 18985 => x"d8a00000", 18986 => x"2b83000c",
    18987 => x"e3ffffe8", 18988 => x"379cfff0", 18989 => x"5b8b0010",
    18990 => x"5b8c000c", 18991 => x"5b8d0008", 18992 => x"5b9d0004",
    18993 => x"b8205800", 18994 => x"44400047", 18995 => x"2822000c",
    18996 => x"58200080", 18997 => x"582000b0", 18998 => x"58220090",
    18999 => x"340c0000", 19000 => x"b9600800", 19001 => x"fbffffaa",
    19002 => x"59610028", 19003 => x"4022003f", 19004 => x"5c400006",
    19005 => x"78040001", 19006 => x"38845ad4", 19007 => x"28230000",
    19008 => x"28820000", 19009 => x"4462005d", 19010 => x"34010000",
    19011 => x"45800030", 19012 => x"3583ffff", 19013 => x"346c0028",
    19014 => x"b58c0800", 19015 => x"b4210800", 19016 => x"b5610800",
    19017 => x"28220000", 19018 => x"5c40000f", 19019 => x"34010000",
    19020 => x"44620027", 19021 => x"34620027", 19022 => x"b4421000",
    19023 => x"b4421000", 19024 => x"b5621000", 19025 => x"e0000002",
    19026 => x"44610044", 19027 => x"28410000", 19028 => x"3463ffff",
    19029 => x"3442fffc", 19030 => x"4420fffc", 19031 => x"596300b0",
    19032 => x"346c0028", 19033 => x"346d0024", 19034 => x"b5ad6800",
    19035 => x"b5ad6800", 19036 => x"b56d6800", 19037 => x"29a20000",
    19038 => x"b9600800", 19039 => x"b58c6000", 19040 => x"fbffff83",
    19041 => x"b58c6000", 19042 => x"b56c1000", 19043 => x"29a40000",
    19044 => x"28430000", 19045 => x"296c00b0", 19046 => x"34840040",
    19047 => x"3463ffff", 19048 => x"59610028", 19049 => x"59a40000",
    19050 => x"58430000", 19051 => x"35830020", 19052 => x"b4631800",
    19053 => x"b4631800", 19054 => x"b5631800", 19055 => x"2824000c",
    19056 => x"28620000", 19057 => x"b4441000", 19058 => x"59620074",
    19059 => x"2b9d0004", 19060 => x"2b8b0010", 19061 => x"2b8c000c",
    19062 => x"2b8d0008", 19063 => x"379c0010", 19064 => x"c3a00000",
    19065 => x"28210028", 19066 => x"296300b0", 19067 => x"34050002",
    19068 => x"4024003f", 19069 => x"eca32800", 19070 => x"64840002",
    19071 => x"a0852000", 19072 => x"4482ffc5", 19073 => x"34620020",
    19074 => x"b4421000", 19075 => x"b4421000", 19076 => x"b5621000",
    19077 => x"28450000", 19078 => x"34640025", 19079 => x"28220004",
    19080 => x"b4842000", 19081 => x"b4842000", 19082 => x"b4a21000",
    19083 => x"b5642000", 19084 => x"58820000", 19085 => x"2824000c",
    19086 => x"34610021", 19087 => x"b4210800", 19088 => x"b4210800",
    19089 => x"b5610800", 19090 => x"b4852800", 19091 => x"346c0001",
    19092 => x"58250000", 19093 => x"e3ffffa3", 19094 => x"34010000",
    19095 => x"596000b0", 19096 => x"2b9d0004", 19097 => x"2b8b0010",
    19098 => x"2b8c000c", 19099 => x"2b8d0008", 19100 => x"379c0010",
    19101 => x"c3a00000", 19102 => x"35820024", 19103 => x"b4421000",
    19104 => x"b4421000", 19105 => x"b5621800", 19106 => x"2c250004",
    19107 => x"28640000", 19108 => x"35820028", 19109 => x"b4421000",
    19110 => x"b4421000", 19111 => x"b5621000", 19112 => x"34a5ffff",
    19113 => x"34840040", 19114 => x"58450000", 19115 => x"58640000",
    19116 => x"596c00b0", 19117 => x"e3ffffbe", 19118 => x"379cffec",
    19119 => x"5b8b0014", 19120 => x"5b8c0010", 19121 => x"5b8d000c",
    19122 => x"5b8e0008", 19123 => x"5b9d0004", 19124 => x"b8406000",
    19125 => x"34020001", 19126 => x"b8205800", 19127 => x"b8607000",
    19128 => x"b8806800", 19129 => x"fbffff73", 19130 => x"b9600800",
    19131 => x"34020000", 19132 => x"fbffff70", 19133 => x"b8202800",
    19134 => x"4420001e", 19135 => x"28a10018", 19136 => x"5c2cfffa",
    19137 => x"28a1001c", 19138 => x"5c2efff8", 19139 => x"28a10020",
    19140 => x"5c2dfff6", 19141 => x"296100b0", 19142 => x"59650028",
    19143 => x"28a2000c", 19144 => x"34210020", 19145 => x"b4210800",
    19146 => x"b4210800", 19147 => x"b5610800", 19148 => x"28230000",
    19149 => x"34010000", 19150 => x"b4431800", 19151 => x"59630074",
    19152 => x"28a30014", 19153 => x"59600078", 19154 => x"34630001",
    19155 => x"c8621000", 19156 => x"59620070", 19157 => x"2b9d0004",
    19158 => x"2b8b0014", 19159 => x"2b8c0010", 19160 => x"2b8d000c",
    19161 => x"2b8e0008", 19162 => x"379c0014", 19163 => x"c3a00000",
    19164 => x"3401fffe", 19165 => x"e3fffff8", 19166 => x"379cfff8",
    19167 => x"5b8b0008", 19168 => x"5b9d0004", 19169 => x"b8205800",
    19170 => x"fbffffcc", 19171 => x"4c200005", 19172 => x"2b9d0004",
    19173 => x"2b8b0008", 19174 => x"379c0008", 19175 => x"c3a00000",
    19176 => x"29610074", 19177 => x"59600028", 19178 => x"2b9d0004",
    19179 => x"2b8b0008", 19180 => x"379c0008", 19181 => x"c3a00000",
    19182 => x"2045ffff", 19183 => x"00460010", 19184 => x"2088ffff",
    19185 => x"00890010", 19186 => x"89053800", 19187 => x"89064000",
    19188 => x"89252800", 19189 => x"00ea0010", 19190 => x"89263000",
    19191 => x"b5052800", 19192 => x"b4aa2800", 19193 => x"50a80003",
    19194 => x"78080001", 19195 => x"b4c83000", 19196 => x"88431000",
    19197 => x"88812000", 19198 => x"00a10010", 19199 => x"3ca50010",
    19200 => x"b4c13000", 19201 => x"20e7ffff", 19202 => x"b4440800",
    19203 => x"b4260800", 19204 => x"b4a71000", 19205 => x"c3a00000",
    19206 => x"44600008", 19207 => x"34040020", 19208 => x"c8832000",
    19209 => x"48800006", 19210 => x"c8041000", 19211 => x"34030000",
    19212 => x"80221000", 19213 => x"b8600800", 19214 => x"c3a00000",
    19215 => x"bc242000", 19216 => x"80431000", 19217 => x"80231800",
    19218 => x"b8821000", 19219 => x"b8600800", 19220 => x"e3fffffa",
    19221 => x"379cfff8", 19222 => x"5b8b0008", 19223 => x"5b9d0004",
    19224 => x"44400022", 19225 => x"b8412000", 19226 => x"3403000f",
    19227 => x"5483000b", 19228 => x"78030001", 19229 => x"38635f4c",
    19230 => x"3c210004", 19231 => x"b4621000", 19232 => x"b4410800",
    19233 => x"40210000", 19234 => x"2b9d0004", 19235 => x"2b8b0008",
    19236 => x"379c0008", 19237 => x"c3a00000", 19238 => x"340b0000",
    19239 => x"4c200003", 19240 => x"c8010800", 19241 => x"340b0001",
    19242 => x"4c400003", 19243 => x"c8021000", 19244 => x"196b0001",
    19245 => x"90c01800", 19246 => x"20630002", 19247 => x"44600008",
    19248 => x"8c220800", 19249 => x"45600002", 19250 => x"c8010800",
    19251 => x"2b9d0004", 19252 => x"2b8b0008", 19253 => x"379c0008",
    19254 => x"c3a00000", 19255 => x"34030000", 19256 => x"f800004a",
    19257 => x"e3fffff8", 19258 => x"90000800", 19259 => x"20210001",
    19260 => x"3c210001", 19261 => x"d0010000", 19262 => x"90e00800",
    19263 => x"bba0f000", 19264 => x"342100a0", 19265 => x"c0200000",
    19266 => x"379cfff8", 19267 => x"5b8b0008", 19268 => x"5b9d0004",
    19269 => x"44400015", 19270 => x"340b0000", 19271 => x"4c200003",
    19272 => x"c8010800", 19273 => x"340b0001", 19274 => x"1443001f",
    19275 => x"90c02000", 19276 => x"98621000", 19277 => x"20840002",
    19278 => x"c8431000", 19279 => x"44800008", 19280 => x"c4220800",
    19281 => x"45600002", 19282 => x"c8010800", 19283 => x"2b9d0004",
    19284 => x"2b8b0008", 19285 => x"379c0008", 19286 => x"c3a00000",
    19287 => x"34030001", 19288 => x"f800002a", 19289 => x"e3fffff8",
    19290 => x"90000800", 19291 => x"20210001", 19292 => x"3c210001",
    19293 => x"d0010000", 19294 => x"90e00800", 19295 => x"bba0f000",
    19296 => x"342100a0", 19297 => x"c0200000", 19298 => x"379cfffc",
    19299 => x"5b9d0004", 19300 => x"44400006", 19301 => x"34030000",
    19302 => x"f800001c", 19303 => x"2b9d0004", 19304 => x"379c0004",
    19305 => x"c3a00000", 19306 => x"90000800", 19307 => x"20210001",
    19308 => x"3c210001", 19309 => x"d0010000", 19310 => x"90e00800",
    19311 => x"bba0f000", 19312 => x"342100a0", 19313 => x"c0200000",
    19314 => x"379cfffc", 19315 => x"5b9d0004", 19316 => x"44400006",
    19317 => x"34030001", 19318 => x"f800000c", 19319 => x"2b9d0004",
    19320 => x"379c0004", 19321 => x"c3a00000", 19322 => x"90000800",
    19323 => x"20210001", 19324 => x"3c210001", 19325 => x"d0010000",
    19326 => x"90e00800", 19327 => x"bba0f000", 19328 => x"342100a0",
    19329 => x"c0200000", 19330 => x"f4222000", 19331 => x"44800018",
    19332 => x"34040001", 19333 => x"4c40000b", 19334 => x"34050000",
    19335 => x"54410003", 19336 => x"c8220800", 19337 => x"b8a42800",
    19338 => x"00840001", 19339 => x"00420001", 19340 => x"5c80fffb",
    19341 => x"5c600002", 19342 => x"b8a00800", 19343 => x"c3a00000",
    19344 => x"3c420001", 19345 => x"3c840001", 19346 => x"f4222800",
    19347 => x"7c860000", 19348 => x"a0c52800", 19349 => x"44a00002",
    19350 => x"4c40fffa", 19351 => x"34050000", 19352 => x"4480fff5",
    19353 => x"34050000", 19354 => x"e3ffffed", 19355 => x"34040001",
    19356 => x"34050000", 19357 => x"e3ffffea", 19358 => x"1422001f",
    19359 => x"98410800", 19360 => x"c8220800", 19361 => x"c3a00000",
    19362 => x"34060003", 19363 => x"b8202000", 19364 => x"b8402800",
    19365 => x"50c3000c", 19366 => x"b8413000", 19367 => x"20c60003",
    19368 => x"5cc0000b", 19369 => x"34010003", 19370 => x"28860000",
    19371 => x"28a20000", 19372 => x"5cc20005", 19373 => x"3463fffc",
    19374 => x"34840004", 19375 => x"34a50004", 19376 => x"5461fffa",
    19377 => x"34010000", 19378 => x"4460000e", 19379 => x"40860000",
    19380 => x"40a10000", 19381 => x"3462ffff", 19382 => x"44c10006",
    19383 => x"e000000a", 19384 => x"40860000", 19385 => x"40a10000",
    19386 => x"3442ffff", 19387 => x"5cc10006", 19388 => x"34840001",
    19389 => x"34a50001", 19390 => x"5c40fffa", 19391 => x"34010000",
    19392 => x"c3a00000", 19393 => x"c8c10800", 19394 => x"c3a00000",
    19395 => x"3404000f", 19396 => x"b8203800", 19397 => x"b8403000",
    19398 => x"5083002d", 19399 => x"b8412000", 19400 => x"20840003",
    19401 => x"5c80002b", 19402 => x"b8402000", 19403 => x"b8202800",
    19404 => x"b8603000", 19405 => x"3407000f", 19406 => x"28880000",
    19407 => x"34c6fff0", 19408 => x"58a80000", 19409 => x"28880004",
    19410 => x"58a80004", 19411 => x"28880008", 19412 => x"58a80008",
    19413 => x"2888000c", 19414 => x"34840010", 19415 => x"58a8000c",
    19416 => x"34a50010", 19417 => x"54c7fff5", 19418 => x"3463fff0",
    19419 => x"00660004", 19420 => x"2063000f", 19421 => x"34c60001",
    19422 => x"3cc60004", 19423 => x"b4263800", 19424 => x"b4463000",
    19425 => x"34020003", 19426 => x"50430011", 19427 => x"34020000",
    19428 => x"34080003", 19429 => x"b4c22000", 19430 => x"28850000",
    19431 => x"b4e22000", 19432 => x"34420004", 19433 => x"58850000",
    19434 => x"c8622000", 19435 => x"5488fffa", 19436 => x"3463fffc",
    19437 => x"00620002", 19438 => x"20630003", 19439 => x"34420001",
    19440 => x"3c420002", 19441 => x"b4e23800", 19442 => x"b4c23000",
    19443 => x"44600008", 19444 => x"34020000", 19445 => x"b4c22000",
    19446 => x"40850000", 19447 => x"b4e22000", 19448 => x"34420001",
    19449 => x"30850000", 19450 => x"5c43fffb", 19451 => x"c3a00000",
    19452 => x"b8203800", 19453 => x"b8403000", 19454 => x"5041000c",
    19455 => x"b4432000", 19456 => x"5024000a", 19457 => x"4460003f",
    19458 => x"b4231000", 19459 => x"3484ffff", 19460 => x"40850000",
    19461 => x"3442ffff", 19462 => x"3463ffff", 19463 => x"30450000",
    19464 => x"5c60fffb", 19465 => x"c3a00000", 19466 => x"3404000f",
    19467 => x"5083002d", 19468 => x"b8412000", 19469 => x"20840003",
    19470 => x"5c80002b", 19471 => x"b8402000", 19472 => x"b8202800",
    19473 => x"b8603000", 19474 => x"3407000f", 19475 => x"28880000",
    19476 => x"34c6fff0", 19477 => x"58a80000", 19478 => x"28880004",
    19479 => x"58a80004", 19480 => x"28880008", 19481 => x"58a80008",
    19482 => x"2888000c", 19483 => x"34840010", 19484 => x"58a8000c",
    19485 => x"34a50010", 19486 => x"54c7fff5", 19487 => x"3463fff0",
    19488 => x"00660004", 19489 => x"2063000f", 19490 => x"34c60001",
    19491 => x"3cc60004", 19492 => x"b4263800", 19493 => x"b4463000",
    19494 => x"34020003", 19495 => x"50430011", 19496 => x"34020000",
    19497 => x"34080003", 19498 => x"b4c22000", 19499 => x"28850000",
    19500 => x"b4e22000", 19501 => x"34420004", 19502 => x"58850000",
    19503 => x"c8622000", 19504 => x"5488fffa", 19505 => x"3463fffc",
    19506 => x"00620002", 19507 => x"20630003", 19508 => x"34420001",
    19509 => x"3c420002", 19510 => x"b4e23800", 19511 => x"b4c23000",
    19512 => x"44600008", 19513 => x"34020000", 19514 => x"b4c22000",
    19515 => x"40850000", 19516 => x"b4e22000", 19517 => x"34420001",
    19518 => x"30850000", 19519 => x"5c43fffb", 19520 => x"c3a00000",
    19521 => x"20250003", 19522 => x"b8202000", 19523 => x"44a0000b",
    19524 => x"4460002c", 19525 => x"3463ffff", 19526 => x"204600ff",
    19527 => x"e0000003", 19528 => x"44600028", 19529 => x"3463ffff",
    19530 => x"30860000", 19531 => x"34840001", 19532 => x"20850003",
    19533 => x"5ca0fffb", 19534 => x"34050003", 19535 => x"50a3001a",
    19536 => x"204500ff", 19537 => x"3ca60008", 19538 => x"340a000f",
    19539 => x"b8c52800", 19540 => x"3ca60010", 19541 => x"b8804000",
    19542 => x"b8c53000", 19543 => x"b8603800", 19544 => x"b8802800",
    19545 => x"3409000f", 19546 => x"546a0017", 19547 => x"34040000",
    19548 => x"34070003", 19549 => x"b5042800", 19550 => x"34840004",
    19551 => x"58a60000", 19552 => x"c8642800", 19553 => x"54a7fffc",
    19554 => x"3463fffc", 19555 => x"00640002", 19556 => x"20630003",
    19557 => x"34840001", 19558 => x"3c840002", 19559 => x"b5044000",
    19560 => x"b9002000", 19561 => x"44600007", 19562 => x"204200ff",
    19563 => x"34050000", 19564 => x"b4853000", 19565 => x"30c20000",
    19566 => x"34a50001", 19567 => x"5c65fffd", 19568 => x"c3a00000",
    19569 => x"58a60000", 19570 => x"58a60004", 19571 => x"58a60008",
    19572 => x"58a6000c", 19573 => x"34e7fff0", 19574 => x"34a50010",
    19575 => x"54e9fffa", 19576 => x"3463fff0", 19577 => x"00680004",
    19578 => x"2063000f", 19579 => x"35080001", 19580 => x"3d080004",
    19581 => x"b4884000", 19582 => x"34040003", 19583 => x"5464ffdc",
    19584 => x"b9002000", 19585 => x"e3ffffe8", 19586 => x"78030001",
    19587 => x"386372b8", 19588 => x"28670000", 19589 => x"b8204800",
    19590 => x"34030000", 19591 => x"34060001", 19592 => x"e0000009",
    19593 => x"40840000", 19594 => x"b4e44000", 19595 => x"41080001",
    19596 => x"21080003", 19597 => x"45060012", 19598 => x"c8a40800",
    19599 => x"5c200013", 19600 => x"44810012", 19601 => x"b5232800",
    19602 => x"40a50000", 19603 => x"b4432000", 19604 => x"34630001",
    19605 => x"b4e54000", 19606 => x"41080001", 19607 => x"21080003",
    19608 => x"5d06fff1", 19609 => x"40840000", 19610 => x"34a50020",
    19611 => x"b4e44000", 19612 => x"41080001", 19613 => x"21080003",
    19614 => x"5d06fff0", 19615 => x"34840020", 19616 => x"c8a40800",
    19617 => x"4420ffef", 19618 => x"c3a00000", 19619 => x"b8411800",
    19620 => x"20630003", 19621 => x"5c60001d", 19622 => x"b8202000",
    19623 => x"28430000", 19624 => x"28210000", 19625 => x"5c230018",
    19626 => x"78030001", 19627 => x"3863604c", 19628 => x"28670000",
    19629 => x"78030001", 19630 => x"38636050", 19631 => x"28660000",
    19632 => x"a4201800", 19633 => x"b4270800", 19634 => x"a0231800",
    19635 => x"a0661800", 19636 => x"34010000", 19637 => x"44600003",
    19638 => x"e000001c", 19639 => x"5c600019", 19640 => x"34840004",
    19641 => x"28810000", 19642 => x"34420004", 19643 => x"28480000",
    19644 => x"b4272800", 19645 => x"a4201800", 19646 => x"a0a31800",
    19647 => x"a0661800", 19648 => x"4428fff7", 19649 => x"b8800800",
    19650 => x"40230000", 19651 => x"5c600006", 19652 => x"e0000009",
    19653 => x"34210001", 19654 => x"40230000", 19655 => x"34420001",
    19656 => x"44600005", 19657 => x"40440000", 19658 => x"4464fffb",
    19659 => x"c8640800", 19660 => x"c3a00000", 19661 => x"40440000",
    19662 => x"c8640800", 19663 => x"c3a00000", 19664 => x"34010000",
    19665 => x"c3a00000", 19666 => x"c3a00000", 19667 => x"b8412800",
    19668 => x"20a50003", 19669 => x"b8403800", 19670 => x"b8202000",
    19671 => x"5ca00018", 19672 => x"78040001", 19673 => x"3884604c",
    19674 => x"28430000", 19675 => x"28880000", 19676 => x"78040001",
    19677 => x"38846050", 19678 => x"28870000", 19679 => x"a4603000",
    19680 => x"b4682000", 19681 => x"a0c43000", 19682 => x"a0c73000",
    19683 => x"b8202000", 19684 => x"5cc5000a", 19685 => x"58830000",
    19686 => x"34420004", 19687 => x"28430000", 19688 => x"34840004",
    19689 => x"a4603000", 19690 => x"b4682800", 19691 => x"a0c52800",
    19692 => x"a0a72800", 19693 => x"44a0fff8", 19694 => x"b8403800",
    19695 => x"34030000", 19696 => x"b4e32800", 19697 => x"40a50000",
    19698 => x"b4833000", 19699 => x"34630001", 19700 => x"30c50000",
    19701 => x"5ca0fffb", 19702 => x"c3a00000", 19703 => x"20220003",
    19704 => x"4440002c", 19705 => x"40230000", 19706 => x"34020000",
    19707 => x"44600027", 19708 => x"b8201000", 19709 => x"e0000003",
    19710 => x"40430000", 19711 => x"44600022", 19712 => x"34420001",
    19713 => x"20430003", 19714 => x"5c60fffc", 19715 => x"78040001",
    19716 => x"3884604c", 19717 => x"28430000", 19718 => x"28860000",
    19719 => x"78040001", 19720 => x"38846050", 19721 => x"28850000",
    19722 => x"a4602000", 19723 => x"b4661800", 19724 => x"a0641800",
    19725 => x"a0651800", 19726 => x"5c600011", 19727 => x"34420004",
    19728 => x"28430000", 19729 => x"b4662000", 19730 => x"a4601800",
    19731 => x"a0831800", 19732 => x"a0651800", 19733 => x"5c60000a",
    19734 => x"34420004", 19735 => x"28430000", 19736 => x"b4662000",
    19737 => x"a4601800", 19738 => x"a0831800", 19739 => x"a0651800",
    19740 => x"4460fff3", 19741 => x"e0000002", 19742 => x"34420001",
    19743 => x"40430000", 19744 => x"5c60fffe", 19745 => x"c8411000",
    19746 => x"b8400800", 19747 => x"c3a00000", 19748 => x"b8201000",
    19749 => x"e3ffffde", 19750 => x"34060000", 19751 => x"44600017",
    19752 => x"b8413800", 19753 => x"20e70003", 19754 => x"3464ffff",
    19755 => x"44e00015", 19756 => x"40230000", 19757 => x"40450000",
    19758 => x"5c65000f", 19759 => x"34060000", 19760 => x"4480000e",
    19761 => x"34210001", 19762 => x"34420001", 19763 => x"5c600004",
    19764 => x"e000000a", 19765 => x"44800033", 19766 => x"44600032",
    19767 => x"40230000", 19768 => x"40450000", 19769 => x"3484ffff",
    19770 => x"34210001", 19771 => x"34420001", 19772 => x"4465fff9",
    19773 => x"c8653000", 19774 => x"b8c00800", 19775 => x"c3a00000",
    19776 => x"b8202800", 19777 => x"34010003", 19778 => x"b8402000",
    19779 => x"50230028", 19780 => x"28a10000", 19781 => x"28420000",
    19782 => x"5c220025", 19783 => x"3463fffc", 19784 => x"b8e03000",
    19785 => x"4460fff5", 19786 => x"78020001", 19787 => x"3842604c",
    19788 => x"28490000", 19789 => x"78020001", 19790 => x"38426050",
    19791 => x"28480000", 19792 => x"a4201000", 19793 => x"b4290800",
    19794 => x"a0220800", 19795 => x"a0280800", 19796 => x"34070003",
    19797 => x"5c20ffe9", 19798 => x"34a50004", 19799 => x"34840004",
    19800 => x"54670006", 19801 => x"b8a00800", 19802 => x"b8801000",
    19803 => x"44600014", 19804 => x"3464ffff", 19805 => x"e3ffffcf",
    19806 => x"28a10000", 19807 => x"288a0000", 19808 => x"b4293000",
    19809 => x"a4201000", 19810 => x"a0c21000", 19811 => x"a0481000",
    19812 => x"5c2a0007", 19813 => x"3463fffc", 19814 => x"44600002",
    19815 => x"4440ffef", 19816 => x"34060000", 19817 => x"b8c00800",
    19818 => x"c3a00000", 19819 => x"b8801000", 19820 => x"b8a00800",
    19821 => x"3464ffff", 19822 => x"e3ffffbe", 19823 => x"40a30000",
    19824 => x"40850000", 19825 => x"c8653000", 19826 => x"e3ffffcc",
    19827 => x"b8412000", 19828 => x"20840003", 19829 => x"74650003",
    19830 => x"64840000", 19831 => x"b8403000", 19832 => x"a0852000",
    19833 => x"b8202800", 19834 => x"44800015", 19835 => x"78040001",
    19836 => x"3884604c", 19837 => x"28890000", 19838 => x"78040001",
    19839 => x"38846050", 19840 => x"28880000", 19841 => x"340a0003",
    19842 => x"e0000006", 19843 => x"58a40000", 19844 => x"3463fffc",
    19845 => x"34a50004", 19846 => x"34420004", 19847 => x"51430007",
    19848 => x"28440000", 19849 => x"a4803800", 19850 => x"b4893000",
    19851 => x"a0e63000", 19852 => x"a0c83000", 19853 => x"44c0fff6",
    19854 => x"b8403000", 19855 => x"44600014", 19856 => x"40c20000",
    19857 => x"3463ffff", 19858 => x"34a40001", 19859 => x"30a20000",
    19860 => x"44400009", 19861 => x"34c20001", 19862 => x"4460000e",
    19863 => x"40450000", 19864 => x"3463ffff", 19865 => x"34420001",
    19866 => x"30850000", 19867 => x"34840001", 19868 => x"5ca0fffa",
    19869 => x"34020000", 19870 => x"44600007", 19871 => x"b4822800",
    19872 => x"30a00000", 19873 => x"34420001", 19874 => x"5c62fffd",
    19875 => x"c3a00000", 19876 => x"c3a00000", 19877 => x"c3a00000",
    19878 => x"34030000", 19879 => x"4440000c", 19880 => x"40240000",
    19881 => x"4480000a", 19882 => x"3442ffff", 19883 => x"b8201800",
    19884 => x"e0000004", 19885 => x"40640000", 19886 => x"3442ffff",
    19887 => x"44800003", 19888 => x"34630001", 19889 => x"5c40fffc",
    19890 => x"c8611800", 19891 => x"b8600800", 19892 => x"c3a00000",
    19893 => x"57522043", 19894 => x"6f72653a", 19895 => x"20737461",
    19896 => x"7274696e", 19897 => x"67207570", 19898 => x"2e2e2e0a",
    19899 => x"00000000", 19900 => x"556e6162", 19901 => x"6c652074",
    19902 => x"6f206465", 19903 => x"7465726d", 19904 => x"696e6520",
    19905 => x"4d414320", 19906 => x"61646472", 19907 => x"6573730a",
    19908 => x"00000000", 19909 => x"4c6f6361", 19910 => x"6c204d41",
    19911 => x"43206164", 19912 => x"64726573", 19913 => x"733a2025",
    19914 => x"3032783a", 19915 => x"25303278", 19916 => x"3a253032",
    19917 => x"783a2530", 19918 => x"32783a25", 19919 => x"3032783a",
    19920 => x"25303278", 19921 => x"0a000000", 19922 => x"73706c6c",
    19923 => x"2d626800", 19924 => x"7368656c", 19925 => x"6c2b6775",
    19926 => x"69000000", 19927 => x"70747000", 19928 => x"75707469",
    19929 => x"6d650000", 19930 => x"63686563", 19931 => x"6b2d6c69",
    19932 => x"6e6b0000", 19933 => x"69646c65", 19934 => x"00000000",
    19935 => x"64696167", 19936 => x"2d66736d", 19937 => x"2d312d25",
    19938 => x"733a2025", 19939 => x"3039642e", 19940 => x"25303364",
    19941 => x"3a200000", 19942 => x"454e5445", 19943 => x"52202573",
    19944 => x"2c207061", 19945 => x"636b6574", 19946 => x"206c656e",
    19947 => x"2025690a", 19948 => x"00000000", 19949 => x"25733a20",
    19950 => x"7265656e", 19951 => x"74657220", 19952 => x"696e2025",
    19953 => x"69206d73", 19954 => x"0a000000", 19955 => x"4c454156",
    19956 => x"45202573", 19957 => x"20286e65", 19958 => x"78743a20",
    19959 => x"25336929", 19960 => x"0a0a0000", 19961 => x"52454356",
    19962 => x"20253032", 19963 => x"64206279", 19964 => x"74657320",
    19965 => x"61742025", 19966 => x"642e2530", 19967 => x"39642028",
    19968 => x"74797065", 19969 => x"2025782c", 19970 => x"20257329",
    19971 => x"0a000000", 19972 => x"66736d20", 19973 => x"666f7220",
    19974 => x"25733a20", 19975 => x"4572726f", 19976 => x"72202569",
    19977 => x"20696e20", 19978 => x"25730a00", 19979 => x"66736d3a",
    19980 => x"20556e6b", 19981 => x"6e6f776e", 19982 => x"20737461",
    19983 => x"74652066", 19984 => x"6f722070", 19985 => x"6f727420",
    19986 => x"25730a00", 19987 => x"70707369", 19988 => x"00000000",
    19989 => x"25732d25", 19990 => x"692d2573", 19991 => x"3a200000",
    19992 => x"25733a20", 19993 => x"6572726f", 19994 => x"72207061",
    19995 => x"7273696e", 19996 => x"67202225", 19997 => x"73220a00",
    19998 => x"64696167", 19999 => x"2d636f6e", 20000 => x"66696700",
    20001 => x"64696167", 20002 => x"2d657874", 20003 => x"656e7369",
    20004 => x"6f6e0000", 20005 => x"64696167", 20006 => x"2d626d63",
    20007 => x"00000000", 20008 => x"64696167", 20009 => x"2d736572",
    20010 => x"766f0000", 20011 => x"64696167", 20012 => x"2d667261",
    20013 => x"6d657300", 20014 => x"64696167", 20015 => x"2d74696d",
    20016 => x"65000000", 20017 => x"64696167", 20018 => x"2d66736d",
    20019 => x"00000000", 20020 => x"50505369", 20021 => x"20666f72",
    20022 => x"20575250", 20023 => x"432e2043", 20024 => x"6f6d6d69",
    20025 => x"74202573", 20026 => x"2c206275", 20027 => x"696c7420",
    20028 => x"6f6e2044", 20029 => x"65632020", 20030 => x"36203230",
    20031 => x"31360a00", 20032 => x"70707369", 20033 => x"2d763230",
    20034 => x"31342e30", 20035 => x"372d3139", 20036 => x"362d6763",
    20037 => x"39336437", 20038 => x"31300000", 20039 => x"50545020",
    20040 => x"73746172", 20041 => x"740a0000", 20042 => x"50545020",
    20043 => x"73746f70", 20044 => x"0a000000", 20045 => x"4c6f636b",
    20046 => x"696e6720", 20047 => x"504c4c00", 20048 => x"0a4c6f63",
    20049 => x"6b207469", 20050 => x"6d656f75", 20051 => x"742e0000",
    20052 => x"2e000000", 20053 => x"77723100", 20054 => x"25732573",
    20055 => x"25303278", 20056 => x"2d253032", 20057 => x"782d2530",
    20058 => x"32782d25", 20059 => x"3032782d", 20060 => x"25303278",
    20061 => x"2d253032", 20062 => x"782d2530", 20063 => x"32782d25",
    20064 => x"3032782d", 20065 => x"25303278", 20066 => x"2d253032",
    20067 => x"780a0000", 20068 => x"25732573", 20069 => x"25732028",
    20070 => x"73697a65", 20071 => x"20256929", 20072 => x"0a000000",
    20073 => x"25732573", 20074 => x"00000000", 20075 => x"25303278",
    20076 => x"00000000", 20077 => x"25735645", 20078 => x"5253494f",
    20079 => x"4e3a2075", 20080 => x"6e737570", 20081 => x"706f7274",
    20082 => x"65642028", 20083 => x"2569290a", 20084 => x"00000000",
    20085 => x"25735645", 20086 => x"5253494f", 20087 => x"4e3a2025",
    20088 => x"69202874", 20089 => x"79706520", 20090 => x"25692c20",
    20091 => x"6c656e20", 20092 => x"25692c20", 20093 => x"646f6d61",
    20094 => x"696e2025", 20095 => x"69290a00", 20096 => x"2573464c",
    20097 => x"4147533a", 20098 => x"20307825", 20099 => x"30347820",
    20100 => x"28636f72", 20101 => x"72656374", 20102 => x"696f6e20",
    20103 => x"2530386c", 20104 => x"75290a00", 20105 => x"504f5254",
    20106 => x"3a200000", 20107 => x"25735245", 20108 => x"53543a20",
    20109 => x"73657120", 20110 => x"25692c20", 20111 => x"6374726c",
    20112 => x"2025692c", 20113 => x"206c6f67", 20114 => x"2d696e74",
    20115 => x"65727661", 20116 => x"6c202569", 20117 => x"0a000000",
    20118 => x"25734d45", 20119 => x"53534147", 20120 => x"453a2028",
    20121 => x"45292053", 20122 => x"594e430a", 20123 => x"00000000",
    20124 => x"25732573", 20125 => x"256c752e", 20126 => x"25303969",
    20127 => x"0a000000", 20128 => x"4d53472d", 20129 => x"53594e43",
    20130 => x"3a200000", 20131 => x"25734d45", 20132 => x"53534147",
    20133 => x"453a2028", 20134 => x"45292044", 20135 => x"454c4159",
    20136 => x"5f524551", 20137 => x"0a000000", 20138 => x"4d53472d",
    20139 => x"44454c41", 20140 => x"595f5245", 20141 => x"513a2000",
    20142 => x"25734d45", 20143 => x"53534147", 20144 => x"453a2028",
    20145 => x"47292046", 20146 => x"4f4c4c4f", 20147 => x"575f5550",
    20148 => x"0a000000", 20149 => x"4d53472d", 20150 => x"464f4c4c",
    20151 => x"4f575f55", 20152 => x"503a2000", 20153 => x"25734d45",
    20154 => x"53534147", 20155 => x"453a2028", 20156 => x"47292044",
    20157 => x"454c4159", 20158 => x"5f524553", 20159 => x"500a0000",
    20160 => x"4d53472d", 20161 => x"44454c41", 20162 => x"595f5245",
    20163 => x"53503a20", 20164 => x"00000000", 20165 => x"25734d45",
    20166 => x"53534147", 20167 => x"453a2028", 20168 => x"47292041",
    20169 => x"4e4e4f55", 20170 => x"4e43450a", 20171 => x"00000000",
    20172 => x"4d53472d", 20173 => x"414e4e4f", 20174 => x"554e4345",
    20175 => x"3a207374", 20176 => x"616d7020", 20177 => x"00000000",
    20178 => x"25732573", 20179 => x"25303278", 20180 => x"2d253032",
    20181 => x"782d2530", 20182 => x"34780a00", 20183 => x"4d53472d",
    20184 => x"414e4e4f", 20185 => x"554e4345", 20186 => x"3a206772",
    20187 => x"616e646d", 20188 => x"61737465", 20189 => x"722d7175",
    20190 => x"616c6974", 20191 => x"79200000", 20192 => x"25734d53",
    20193 => x"472d414e", 20194 => x"4e4f554e", 20195 => x"43453a20",
    20196 => x"6772616e", 20197 => x"646d6173", 20198 => x"7465722d",
    20199 => x"7072696f", 20200 => x"20256920", 20201 => x"25690a00",
    20202 => x"25732573", 20203 => x"25303278", 20204 => x"2d253032",
    20205 => x"782d2530", 20206 => x"32782d25", 20207 => x"3032782d",
    20208 => x"25303278", 20209 => x"2d253032", 20210 => x"782d2530",
    20211 => x"32782d25", 20212 => x"3032780a", 20213 => x"00000000",
    20214 => x"4d53472d", 20215 => x"414e4e4f", 20216 => x"554e4345",
    20217 => x"3a206772", 20218 => x"616e646d", 20219 => x"61737465",
    20220 => x"722d6964", 20221 => x"20000000", 20222 => x"25734d45",
    20223 => x"53534147", 20224 => x"453a2028", 20225 => x"47292053",
    20226 => x"49474e41", 20227 => x"4c494e47", 20228 => x"0a000000",
    20229 => x"4d53472d", 20230 => x"5349474e", 20231 => x"414c494e",
    20232 => x"473a2074", 20233 => x"61726765", 20234 => x"742d706f",
    20235 => x"72742000", 20236 => x"2573544c", 20237 => x"563a2074",
    20238 => x"6f6f2073", 20239 => x"686f7274", 20240 => x"20282569",
    20241 => x"202d2025", 20242 => x"69203d20", 20243 => x"2569290a",
    20244 => x"00000000", 20245 => x"2573544c", 20246 => x"563a2074",
    20247 => x"79706520", 20248 => x"25303478", 20249 => x"206c656e",
    20250 => x"20256920", 20251 => x"6f756920", 20252 => x"25303278",
    20253 => x"3a253032", 20254 => x"783a2530", 20255 => x"32782073",
    20256 => x"75622025", 20257 => x"3032783a", 20258 => x"25303278",
    20259 => x"3a253032", 20260 => x"780a0000", 20261 => x"2573544c",
    20262 => x"563a2074", 20263 => x"6f6f2073", 20264 => x"686f7274",
    20265 => x"20286578", 20266 => x"70656374", 20267 => x"65642025",
    20268 => x"692c2074", 20269 => x"6f74616c", 20270 => x"20256929",
    20271 => x"0a000000", 20272 => x"544c563a", 20273 => x"20000000",
    20274 => x"746c762d", 20275 => x"636f6e74", 20276 => x"656e7400",
    20277 => x"44554d50", 20278 => x"3a200000", 20279 => x"7061796c",
    20280 => x"6f616400", 20281 => x"20696e76", 20282 => x"616c6964",
    20283 => x"00000000", 20284 => x"25735449", 20285 => x"4d453a20",
    20286 => x"28256c69", 20287 => x"202d2030", 20288 => x"78256c78",
    20289 => x"2920256c", 20290 => x"692e2530", 20291 => x"366c6925",
    20292 => x"730a0000", 20293 => x"2573564c", 20294 => x"414e2025",
    20295 => x"690a0000", 20296 => x"25734554", 20297 => x"483a2025",
    20298 => x"30347820", 20299 => x"28253032", 20300 => x"783a2530",
    20301 => x"32783a25", 20302 => x"3032783a", 20303 => x"25303278",
    20304 => x"3a253032", 20305 => x"783a2530", 20306 => x"3278202d",
    20307 => x"3e202530", 20308 => x"32783a25", 20309 => x"3032783a",
    20310 => x"25303278", 20311 => x"3a253032", 20312 => x"783a2530",
    20313 => x"32783a25", 20314 => x"30327829", 20315 => x"0a000000",
    20316 => x"25734950", 20317 => x"3a202569", 20318 => x"20282569",
    20319 => x"2e25692e", 20320 => x"25692e25", 20321 => x"69202d3e",
    20322 => x"2025692e", 20323 => x"25692e25", 20324 => x"692e2569",
    20325 => x"29206c65", 20326 => x"6e202569", 20327 => x"0a000000",
    20328 => x"25735544", 20329 => x"503a2028", 20330 => x"2569202d",
    20331 => x"3e202569", 20332 => x"29206c65", 20333 => x"6e202569",
    20334 => x"0a000000", 20335 => x"25733a20", 20336 => x"256c690a",
    20337 => x"00000000", 20338 => x"5761726e", 20339 => x"696e673a",
    20340 => x"2025733a", 20341 => x"2063616e", 20342 => x"206e6f74",
    20343 => x"2061646a", 20344 => x"75737420", 20345 => x"66726571",
    20346 => x"5f707062", 20347 => x"20256c69", 20348 => x"0a000000",
    20349 => x"25733a20", 20350 => x"25396c75", 20351 => x"2e253039",
    20352 => x"6c690a00", 20353 => x"25733a20", 20354 => x"736e743d",
    20355 => x"25642c20", 20356 => x"7365633d", 20357 => x"25642c20",
    20358 => x"6e736563", 20359 => x"3d25640a", 20360 => x"00000000",
    20361 => x"73656e64", 20362 => x"3a200000", 20363 => x"72656376",
    20364 => x"3a200000", 20365 => x"696e6974", 20366 => x"69616c69",
    20367 => x"7a696e67", 20368 => x"00000000", 20369 => x"6661756c",
    20370 => x"74790000", 20371 => x"64697361", 20372 => x"626c6564",
    20373 => x"00000000", 20374 => x"6c697374", 20375 => x"656e696e",
    20376 => x"67000000", 20377 => x"756e6361", 20378 => x"6c696272",
    20379 => x"61746564", 20380 => x"00000000", 20381 => x"736c6176",
    20382 => x"65000000", 20383 => x"756e6361", 20384 => x"6c696272",
    20385 => x"61746564", 20386 => x"2f77722d", 20387 => x"70726573",
    20388 => x"656e7400", 20389 => x"6d617374", 20390 => x"65722f77",
    20391 => x"722d6d2d", 20392 => x"6c6f636b", 20393 => x"00000000",
    20394 => x"756e6361", 20395 => x"6c696272", 20396 => x"61746564",
    20397 => x"2f77722d", 20398 => x"732d6c6f", 20399 => x"636b0000",
    20400 => x"756e6361", 20401 => x"6c696272", 20402 => x"61746564",
    20403 => x"2f77722d", 20404 => x"6c6f636b", 20405 => x"65640000",
    20406 => x"77722d63", 20407 => x"616c6962", 20408 => x"72617469",
    20409 => x"6f6e0000", 20410 => x"77722d63", 20411 => x"616c6962",
    20412 => x"72617465", 20413 => x"64000000", 20414 => x"77722d72",
    20415 => x"6573702d", 20416 => x"63616c69", 20417 => x"622d7265",
    20418 => x"71000000", 20419 => x"77722d6c", 20420 => x"696e6b2d",
    20421 => x"6f6e0000", 20422 => x"686f6f6b", 20423 => x"3a202573",
    20424 => x"0a000000", 20425 => x"5432206f", 20426 => x"72205433",
    20427 => x"20696e63", 20428 => x"6f727265", 20429 => x"63742c20",
    20430 => x"64697363", 20431 => x"61726469", 20432 => x"6e672074",
    20433 => x"75706c65", 20434 => x"0a000000", 20435 => x"48616e64",
    20436 => x"7368616b", 20437 => x"65206661", 20438 => x"696c7572",
    20439 => x"653a206e", 20440 => x"6f77206e", 20441 => x"6f6e2d77",
    20442 => x"72202573", 20443 => x"0a000000", 20444 => x"52657472",
    20445 => x"79206f6e", 20446 => x"2074696d", 20447 => x"656f7574",
    20448 => x"0a000000", 20449 => x"25733a20", 20450 => x"73756273",
    20451 => x"74617465", 20452 => x"2025690a", 20453 => x"00000000",
    20454 => x"54783d3e", 20455 => x"3e736361", 20456 => x"6c656450",
    20457 => x"69636f73", 20458 => x"65636f6e", 20459 => x"64732e6d",
    20460 => x"7362203d", 20461 => x"20307825", 20462 => x"780a0000",
    20463 => x"54783d3e", 20464 => x"3e736361", 20465 => x"6c656450",
    20466 => x"69636f73", 20467 => x"65636f6e", 20468 => x"64732e6c",
    20469 => x"7362203d", 20470 => x"20307825", 20471 => x"780a0000",
    20472 => x"52782066", 20473 => x"69786564", 20474 => x"2064656c",
    20475 => x"6179203d", 20476 => x"2025640a", 20477 => x"00000000",
    20478 => x"52783d3e", 20479 => x"3e736361", 20480 => x"6c656450",
    20481 => x"69636f73", 20482 => x"65636f6e", 20483 => x"64732e6d",
    20484 => x"7362203d", 20485 => x"20307825", 20486 => x"780a0000",
    20487 => x"52783d3e", 20488 => x"3e736361", 20489 => x"6c656450",
    20490 => x"69636f73", 20491 => x"65636f6e", 20492 => x"64732e6c",
    20493 => x"7362203d", 20494 => x"20307825", 20495 => x"780a0000",
    20496 => x"4552524f", 20497 => x"523a204e", 20498 => x"65772063",
    20499 => x"6c617373", 20500 => x"2025690a", 20501 => x"00000000",
    20502 => x"4255473a", 20503 => x"20547279", 20504 => x"696e6720",
    20505 => x"746f2073", 20506 => x"656e6420", 20507 => x"696e7661",
    20508 => x"6c696420", 20509 => x"77725f6d", 20510 => x"7367206d",
    20511 => x"6f64653d", 20512 => x"25782069", 20513 => x"643d2578",
    20514 => x"00000000", 20515 => x"68616e64", 20516 => x"6c652053",
    20517 => x"69676e61", 20518 => x"6c696e67", 20519 => x"206d7367",
    20520 => x"2c206661", 20521 => x"696c6564", 20522 => x"2c205468",
    20523 => x"69732069", 20524 => x"73206e6f", 20525 => x"74206f72",
    20526 => x"67616e69", 20527 => x"7a617469", 20528 => x"6f6e2065",
    20529 => x"7874656e", 20530 => x"73696f6e", 20531 => x"20544c56",
    20532 => x"203d2030", 20533 => x"7825780a", 20534 => x"00000000",
    20535 => x"68616e64", 20536 => x"6c652053", 20537 => x"69676e61",
    20538 => x"6c696e67", 20539 => x"206d7367", 20540 => x"2c206661",
    20541 => x"696c6564", 20542 => x"2c206e6f", 20543 => x"74204345",
    20544 => x"524e2773", 20545 => x"204f5549", 20546 => x"203d2030",
    20547 => x"7825780a", 20548 => x"00000000", 20549 => x"68616e64",
    20550 => x"6c652053", 20551 => x"69676e61", 20552 => x"6c696e67",
    20553 => x"206d7367", 20554 => x"2c206661", 20555 => x"696c6564",
    20556 => x"2c206e6f", 20557 => x"74205768", 20558 => x"69746520",
    20559 => x"52616262", 20560 => x"6974206d", 20561 => x"61676963",
    20562 => x"206e756d", 20563 => x"62657220", 20564 => x"3d203078",
    20565 => x"25780a00", 20566 => x"68616e64", 20567 => x"6c652053",
    20568 => x"69676e61", 20569 => x"6c696e67", 20570 => x"206d7367",
    20571 => x"2c206661", 20572 => x"696c6564", 20573 => x"2c206e6f",
    20574 => x"74207375", 20575 => x"70706f72", 20576 => x"74656420",
    20577 => x"76657273", 20578 => x"696f6e20", 20579 => x"6e756d62",
    20580 => x"6572203d", 20581 => x"20307825", 20582 => x"780a0000",
    20583 => x"25732825", 20584 => x"6429204d", 20585 => x"65737361",
    20586 => x"67652063", 20587 => x"616e2774", 20588 => x"20626520",
    20589 => x"73656e74", 20590 => x"0a000000", 20591 => x"53454e54",
    20592 => x"20253032", 20593 => x"64206279", 20594 => x"74657320",
    20595 => x"61742025", 20596 => x"642e2530", 20597 => x"39642028",
    20598 => x"2573290a", 20599 => x"00000000", 20600 => x"556e696e",
    20601 => x"69746961", 20602 => x"6c697a65", 20603 => x"64000000",
    20604 => x"20287761", 20605 => x"69742066", 20606 => x"6f722068",
    20607 => x"77290000", 20608 => x"4552524f", 20609 => x"523a2025",
    20610 => x"733a2054", 20611 => x"696d6573", 20612 => x"74616d70",
    20613 => x"73496e63", 20614 => x"6f727265", 20615 => x"63743a20",
    20616 => x"25642025", 20617 => x"64202564", 20618 => x"2025640a",
    20619 => x"00000000", 20620 => x"2573203d", 20621 => x"2025643a",
    20622 => x"25643a25", 20623 => x"640a0000", 20624 => x"73657276",
    20625 => x"6f3a7431", 20626 => x"00000000", 20627 => x"73657276",
    20628 => x"6f3a7432", 20629 => x"00000000", 20630 => x"73657276",
    20631 => x"6f3a7433", 20632 => x"00000000", 20633 => x"73657276",
    20634 => x"6f3a7434", 20635 => x"00000000", 20636 => x"2d3e6d64",
    20637 => x"656c6179", 20638 => x"00000000", 20639 => x"504c4c20",
    20640 => x"4f75744f", 20641 => x"664c6f63", 20642 => x"6b2c2073",
    20643 => x"686f756c", 20644 => x"64207265", 20645 => x"73746172",
    20646 => x"74207379", 20647 => x"6e630a00", 20648 => x"73657276",
    20649 => x"6f3a6275", 20650 => x"73790a00", 20651 => x"6f666673",
    20652 => x"65745f68", 20653 => x"773a2025", 20654 => x"6c692e25",
    20655 => x"30396c69", 20656 => x"20282b25", 20657 => x"6c69290a",
    20658 => x"00000000", 20659 => x"77725f73", 20660 => x"6572766f",
    20661 => x"20737461", 20662 => x"74653a20", 20663 => x"25732573",
    20664 => x"0a000000", 20665 => x"6f6c6473", 20666 => x"65747020",
    20667 => x"25692c20", 20668 => x"6f666673", 20669 => x"65742025",
    20670 => x"693a2530", 20671 => x"34690a00", 20672 => x"61646a75",
    20673 => x"73742070", 20674 => x"68617365", 20675 => x"2025690a",
    20676 => x"00000000", 20677 => x"53594e43", 20678 => x"5f4e5345",
    20679 => x"43000000", 20680 => x"53594e43", 20681 => x"5f534543",
    20682 => x"00000000", 20683 => x"53594e43", 20684 => x"5f504841",
    20685 => x"53450000", 20686 => x"54524143", 20687 => x"4b5f5048",
    20688 => x"41534500", 20689 => x"57414954", 20690 => x"5f4f4646",
    20691 => x"5345545f", 20692 => x"53544142", 20693 => x"4c450000",
    20694 => x"7072652d", 20695 => x"6d617374", 20696 => x"65720000",
    20697 => x"70617373", 20698 => x"69766500", 20699 => x"25733a20",
    20700 => x"63616e27", 20701 => x"7420696e", 20702 => x"69742065",
    20703 => x"7874656e", 20704 => x"73696f6e", 20705 => x"0a000000",
    20706 => x"636c6f63", 20707 => x"6b20636c", 20708 => x"61737320",
    20709 => x"3d202564", 20710 => x"0a000000", 20711 => x"636c6f63",
    20712 => x"6b206163", 20713 => x"63757261", 20714 => x"6379203d",
    20715 => x"2025640a", 20716 => x"00000000", 20717 => x"70705f73",
    20718 => x"6c617665", 20719 => x"203a2044", 20720 => x"656c6179",
    20721 => x"20526573", 20722 => x"7020646f", 20723 => x"65736e27",
    20724 => x"74206d61", 20725 => x"74636820", 20726 => x"44656c61",
    20727 => x"79205265", 20728 => x"710a0000", 20729 => x"4e657720",
    20730 => x"666f7265", 20731 => x"69676e20", 20732 => x"4d617374",
    20733 => x"65722025", 20734 => x"69206164", 20735 => x"6465640a",
    20736 => x"00000000", 20737 => x"4552524f", 20738 => x"523a2025",
    20739 => x"733a2046", 20740 => x"6f6c6c6f", 20741 => x"77207570",
    20742 => x"206d6573", 20743 => x"73616765", 20744 => x"20697320",
    20745 => x"6e6f7420", 20746 => x"66726f6d", 20747 => x"20637572",
    20748 => x"72656e74", 20749 => x"20706172", 20750 => x"656e740a",
    20751 => x"00000000", 20752 => x"4552524f", 20753 => x"523a2025",
    20754 => x"733a2053", 20755 => x"6c617665", 20756 => x"20776173",
    20757 => x"206e6f74", 20758 => x"20776169", 20759 => x"74696e67",
    20760 => x"20612066", 20761 => x"6f6c6c6f", 20762 => x"77207570",
    20763 => x"206d6573", 20764 => x"73616765", 20765 => x"0a000000",
    20766 => x"4552524f", 20767 => x"523a2025", 20768 => x"733a2053",
    20769 => x"65717565", 20770 => x"6e636549", 20771 => x"44202564",
    20772 => x"20646f65", 20773 => x"736e2774", 20774 => x"206d6174",
    20775 => x"6368206c", 20776 => x"61737420", 20777 => x"53796e63",
    20778 => x"206d6573", 20779 => x"73616765", 20780 => x"2025640a",
    20781 => x"00000000", 20782 => x"416e6e6f", 20783 => x"756e6365",
    20784 => x"206d6573", 20785 => x"73616765", 20786 => x"2066726f",
    20787 => x"6d20616e", 20788 => x"6f746865", 20789 => x"7220666f",
    20790 => x"72656967", 20791 => x"6e206d61", 20792 => x"73746572",
    20793 => x"0a000000", 20794 => x"25733a25", 20795 => x"693a2045",
    20796 => x"72726f72", 20797 => x"20310a00", 20798 => x"25733a25",
    20799 => x"693a2045", 20800 => x"72726f72", 20801 => x"20320a00",
    20802 => x"42657374", 20803 => x"20666f72", 20804 => x"6569676e",
    20805 => x"206d6173", 20806 => x"74657220", 20807 => x"69732025",
    20808 => x"692f2569", 20809 => x"0a000000", 20810 => x"25733a20",
    20811 => x"6572726f", 20812 => x"720a0000", 20813 => x"25733a20",
    20814 => x"70617373", 20815 => x"6976650a", 20816 => x"00000000",
    20817 => x"25733a20", 20818 => x"6d617374", 20819 => x"65720a00",
    20820 => x"4e657720", 20821 => x"55544320", 20822 => x"6f666673",
    20823 => x"65743a20", 20824 => x"25690a00", 20825 => x"25733a20",
    20826 => x"736c6176", 20827 => x"650a0000", 20828 => x"73796e63",
    20829 => x"00000000", 20830 => x"64656c61", 20831 => x"795f7265",
    20832 => x"71000000", 20833 => x"7064656c", 20834 => x"61795f72",
    20835 => x"65710000", 20836 => x"7064656c", 20837 => x"61795f72",
    20838 => x"65737000", 20839 => x"64656c61", 20840 => x"795f7265",
    20841 => x"73700000", 20842 => x"7064656c", 20843 => x"61795f72",
    20844 => x"6573705f", 20845 => x"666f6c6c", 20846 => x"6f775f75",
    20847 => x"70000000", 20848 => x"616e6e6f", 20849 => x"756e6365",
    20850 => x"00000000", 20851 => x"7369676e", 20852 => x"616c696e",
    20853 => x"67000000", 20854 => x"6d616e61", 20855 => x"67656d65",
    20856 => x"6e740000", 20857 => x"4552524f", 20858 => x"523a2042",
    20859 => x"55473a20", 20860 => x"25732064", 20861 => x"6f65736e",
    20862 => x"27742073", 20863 => x"7570706f", 20864 => x"7274206e",
    20865 => x"65676174", 20866 => x"69766573", 20867 => x"0a000000",
    20868 => x"4552524f", 20869 => x"523a204e", 20870 => x"65676174",
    20871 => x"69766520", 20872 => x"76616c75", 20873 => x"65206361",
    20874 => x"6e6e6f74", 20875 => x"20626520", 20876 => x"636f6e76",
    20877 => x"65727465", 20878 => x"6420696e", 20879 => x"746f2074",
    20880 => x"696d6573", 20881 => x"74616d70", 20882 => x"0a000000",
    20883 => x"4552524f", 20884 => x"523a2074", 20885 => x"6f5f5469",
    20886 => x"6d65496e", 20887 => x"7465726e", 20888 => x"616c3a20",
    20889 => x"7365636f", 20890 => x"6e647320", 20891 => x"6669656c",
    20892 => x"64206973", 20893 => x"20686967", 20894 => x"68657220",
    20895 => x"7468616e", 20896 => x"20736967", 20897 => x"6e656420",
    20898 => x"696e7465", 20899 => x"67657220", 20900 => x"28333262",
    20901 => x"69747329", 20902 => x"0a000000", 20903 => x"2d000000",
    20904 => x"25732564", 20905 => x"2e253039", 20906 => x"64000000",
    20907 => x"6572726f", 20908 => x"7220696e", 20909 => x"20745f6f",
    20910 => x"70732d3e", 20911 => x"73657276", 20912 => x"6f5f696e",
    20913 => x"69740000", 20914 => x"496e6974", 20915 => x"69616c69",
    20916 => x"7a65643a", 20917 => x"206f6273", 20918 => x"5f647269",
    20919 => x"66742025", 20920 => x"6c6c690a", 20921 => x"00000000",
    20922 => x"636f7272", 20923 => x"65637469", 20924 => x"6f6e2066",
    20925 => x"69656c64", 20926 => x"20313a20", 20927 => x"25730a00",
    20928 => x"64697363", 20929 => x"61726420", 20930 => x"54332f54",
    20931 => x"343a2077", 20932 => x"65206d69", 20933 => x"73732054",
    20934 => x"312f5432", 20935 => x"0a000000", 20936 => x"636f7272",
    20937 => x"65637469", 20938 => x"6f6e2066", 20939 => x"69656c64",
    20940 => x"20323a20", 20941 => x"25730a00", 20942 => x"54313a20",
    20943 => x"25730a00", 20944 => x"54323a20", 20945 => x"25730a00",
    20946 => x"54333a20", 20947 => x"25730a00", 20948 => x"54343a20",
    20949 => x"25730a00", 20950 => x"4d617374", 20951 => x"65722074",
    20952 => x"6f20736c", 20953 => x"6176653a", 20954 => x"2025730a",
    20955 => x"00000000", 20956 => x"536c6176", 20957 => x"6520746f",
    20958 => x"206d6173", 20959 => x"7465723a", 20960 => x"2025730a",
    20961 => x"00000000", 20962 => x"6d65616e", 20963 => x"50617468",
    20964 => x"44656c61", 20965 => x"793a2025", 20966 => x"730a0000",
    20967 => x"73657276", 20968 => x"6f206162", 20969 => x"6f727465",
    20970 => x"642c2064", 20971 => x"656c6179", 20972 => x"20677265",
    20973 => x"61746572", 20974 => x"20746861", 20975 => x"6e203120",
    20976 => x"7365636f", 20977 => x"6e640a00", 20978 => x"73657276",
    20979 => x"6f206162", 20980 => x"6f727465", 20981 => x"642c2064",
    20982 => x"656c6179", 20983 => x"20256420", 20984 => x"6f722025",
    20985 => x"64206772", 20986 => x"65617465", 20987 => x"72207468",
    20988 => x"616e2063", 20989 => x"6f6e6669", 20990 => x"67757265",
    20991 => x"64206d61", 20992 => x"78696d75", 20993 => x"6d202564",
    20994 => x"0a000000", 20995 => x"5472696d", 20996 => x"20746f6f",
    20997 => x"2d6c6f6e", 20998 => x"67206d70", 20999 => x"643a2025",
    21000 => x"690a0000", 21001 => x"41667465", 21002 => x"72206176",
    21003 => x"67282569", 21004 => x"292c206d", 21005 => x"65616e50",
    21006 => x"61746844", 21007 => x"656c6179", 21008 => x"3a202569",
    21009 => x"0a000000", 21010 => x"4f666673", 21011 => x"65742066",
    21012 => x"726f6d20", 21013 => x"6d617374", 21014 => x"65723a20",
    21015 => x"20202020", 21016 => x"25730a00", 21017 => x"73657276",
    21018 => x"6f206162", 21019 => x"6f727465", 21020 => x"642c206f",
    21021 => x"66667365", 21022 => x"74206772", 21023 => x"65617465",
    21024 => x"72207468", 21025 => x"616e2031", 21026 => x"20736563",
    21027 => x"6f6e640a", 21028 => x"00000000", 21029 => x"73657276",
    21030 => x"6f206162", 21031 => x"6f727465", 21032 => x"642c206f",
    21033 => x"66667365", 21034 => x"74206772", 21035 => x"65617465",
    21036 => x"72207468", 21037 => x"616e2063", 21038 => x"6f6e6669",
    21039 => x"67757265", 21040 => x"64206d61", 21041 => x"78696d75",
    21042 => x"6d202564", 21043 => x"0a000000", 21044 => x"4f627365",
    21045 => x"72766564", 21046 => x"20647269", 21047 => x"66743a20",
    21048 => x"2539690a", 21049 => x"00000000", 21050 => x"74696d65",
    21051 => x"6f757420", 21052 => x"65787069", 21053 => x"7265643a",
    21054 => x"2025730a", 21055 => x"00000000", 21056 => x"50505f54",
    21057 => x"4f5f4445", 21058 => x"4c415952", 21059 => x"45510000",
    21060 => x"50505f54", 21061 => x"4f5f5359", 21062 => x"4e430000",
    21063 => x"50505f54", 21064 => x"4f5f414e", 21065 => x"4e5f5245",
    21066 => x"43454950", 21067 => x"54000000", 21068 => x"50505f54",
    21069 => x"4f5f414e", 21070 => x"4e5f494e", 21071 => x"54455256",
    21072 => x"414c0000", 21073 => x"50505f54", 21074 => x"4f5f4641",
    21075 => x"554c5459", 21076 => x"00000000", 21077 => x"50505f54",
    21078 => x"4f5f4558", 21079 => x"545f3000", 21080 => x"50505f54",
    21081 => x"4f5f4558", 21082 => x"545f3100", 21083 => x"50505f54",
    21084 => x"4f5f4558", 21085 => x"545f3200", 21086 => x"536c6176",
    21087 => x"65204f6e", 21088 => x"6c792c20", 21089 => x"636c6f63",
    21090 => x"6b20636c", 21091 => x"61737320", 21092 => x"73657420",
    21093 => x"746f2032", 21094 => x"35350a00", 21095 => x"25750000",
    21096 => x"25752575", 21097 => x"00000000", 21098 => x"6c6e6b3a",
    21099 => x"25642072", 21100 => x"783a2564", 21101 => x"2074783a",
    21102 => x"25642000", 21103 => x"6c6f636b", 21104 => x"3a256420",
    21105 => x"00000000", 21106 => x"7074703a", 21107 => x"25732000",
    21108 => x"73763a25", 21109 => x"64200000", 21110 => x"73733a27",
    21111 => x"25732720", 21112 => x"00000000", 21113 => x"6175783a",
    21114 => x"25782000", 21115 => x"7365633a", 21116 => x"2564206e",
    21117 => x"7365633a", 21118 => x"25642000", 21119 => x"6d753a25",
    21120 => x"73200000", 21121 => x"646d733a", 21122 => x"25732000",
    21123 => x"6474786d", 21124 => x"3a256420", 21125 => x"6472786d",
    21126 => x"3a256420", 21127 => x"00000000", 21128 => x"64747873",
    21129 => x"3a256420", 21130 => x"64727873", 21131 => x"3a256420",
    21132 => x"00000000", 21133 => x"6173796d", 21134 => x"3a256420",
    21135 => x"00000000", 21136 => x"63727474", 21137 => x"3a257320",
    21138 => x"00000000", 21139 => x"636b6f3a", 21140 => x"25642000",
    21141 => x"73657470", 21142 => x"3a256420", 21143 => x"00000000",
    21144 => x"75636e74", 21145 => x"3a256420", 21146 => x"00000000",
    21147 => x"68643a25", 21148 => x"64206d64", 21149 => x"3a256420",
    21150 => x"61643a25", 21151 => x"64200000", 21152 => x"70636200",
    21153 => x"74656d70", 21154 => x"3a202564", 21155 => x"2e253034",
    21156 => x"64204300", 21157 => x"0a0a5054", 21158 => x"50207374",
    21159 => x"61747573", 21160 => x"3a200000", 21161 => x"25730000",
    21162 => x"0a0a5379", 21163 => x"6e632069", 21164 => x"6e666f20",
    21165 => x"6e6f7420", 21166 => x"76616c69", 21167 => x"640a0a00",
    21168 => x"0a0a5379", 21169 => x"6e636872", 21170 => x"6f6e697a",
    21171 => x"6174696f", 21172 => x"6e207374", 21173 => x"61747573",
    21174 => x"3a0a0a00", 21175 => x"57522050", 21176 => x"54502043",
    21177 => x"6f726520", 21178 => x"53796e63", 21179 => x"204d6f6e",
    21180 => x"69746f72", 21181 => x"20762031", 21182 => x"2e300000",
    21183 => x"45736320", 21184 => x"3d206578", 21185 => x"69740000",
    21186 => x"0a0a5441", 21187 => x"49205469", 21188 => x"6d653a20",
    21189 => x"20202020", 21190 => x"20202020", 21191 => x"20202020",
    21192 => x"20202020", 21193 => x"20000000", 21194 => x"0a0a4c69",
    21195 => x"6e6b2073", 21196 => x"74617475", 21197 => x"733a0000",
    21198 => x"25733a20", 21199 => x"00000000", 21200 => x"77727531",
    21201 => x"00000000", 21202 => x"4c696e6b", 21203 => x"20757020",
    21204 => x"20200000", 21205 => x"4c696e6b", 21206 => x"20646f77",
    21207 => x"6e200000", 21208 => x"2852583a", 21209 => x"2025642c",
    21210 => x"2054583a", 21211 => x"20256429", 21212 => x"2c206d6f",
    21213 => x"64653a20", 21214 => x"00000000", 21215 => x"5752204f",
    21216 => x"66660000", 21217 => x"436c6f63", 21218 => x"6b206f66",
    21219 => x"66736574", 21220 => x"3a202020", 21221 => x"20202020",
    21222 => x"20202020", 21223 => x"20202020", 21224 => x"20200000",
    21225 => x"2532692e", 21226 => x"25303969", 21227 => x"20730000",
    21228 => x"25396920", 21229 => x"6e730000", 21230 => x"0a4f6e65",
    21231 => x"2d776179", 21232 => x"2064656c", 21233 => x"61792061",
    21234 => x"76657261", 21235 => x"6765643a", 21236 => x"20202020",
    21237 => x"20202000", 21238 => x"0a4f6273", 21239 => x"65727665",
    21240 => x"64206472", 21241 => x"6966743a", 21242 => x"20202020",
    21243 => x"20202020", 21244 => x"20202020", 21245 => x"20202000",
    21246 => x"5752204d", 21247 => x"61737465", 21248 => x"72202000",
    21249 => x"57522053", 21250 => x"6c617665", 21251 => x"20202000",
    21252 => x"57522055", 21253 => x"6e6b6e6f", 21254 => x"776e2020",
    21255 => x"20000000", 21256 => x"4c6f636b", 21257 => x"65642020",
    21258 => x"00000000", 21259 => x"4e6f4c6f", 21260 => x"636b2020",
    21261 => x"00000000", 21262 => x"43616c69", 21263 => x"62726174",
    21264 => x"65642020", 21265 => x"00000000", 21266 => x"556e6361",
    21267 => x"6c696272", 21268 => x"61746564", 21269 => x"20200000",
    21270 => x"0a495076", 21271 => x"343a2000", 21272 => x"424f4f54",
    21273 => x"50207275", 21274 => x"6e6e696e", 21275 => x"67000000",
    21276 => x"25732028", 21277 => x"66726f6d", 21278 => x"20626f6f",
    21279 => x"74702900", 21280 => x"25732028", 21281 => x"73746174",
    21282 => x"69632061", 21283 => x"73736967", 21284 => x"6e6d656e",
    21285 => x"74290000", 21286 => x"53657276", 21287 => x"6f207374",
    21288 => x"6174653a", 21289 => x"20202020", 21290 => x"20202020",
    21291 => x"20202020", 21292 => x"20202000", 21293 => x"50686173",
    21294 => x"65207472", 21295 => x"61636b69", 21296 => x"6e673a20",
    21297 => x"20202020", 21298 => x"20202020", 21299 => x"20202000",
    21300 => x"4f4e0a00", 21301 => x"4f46460a", 21302 => x"00000000",
    21303 => x"41757820", 21304 => x"636c6f63", 21305 => x"6b207374",
    21306 => x"61747573", 21307 => x"3a202020", 21308 => x"20202020",
    21309 => x"20202000", 21310 => x"656e6162", 21311 => x"6c656400",
    21312 => x"2c206c6f", 21313 => x"636b6564", 21314 => x"00000000",
    21315 => x"0a54696d", 21316 => x"696e6720", 21317 => x"70617261",
    21318 => x"6d657465", 21319 => x"72733a0a", 21320 => x"0a000000",
    21321 => x"526f756e", 21322 => x"642d7472", 21323 => x"69702074",
    21324 => x"696d6520", 21325 => x"286d7529", 21326 => x"3a202020",
    21327 => x"20000000", 21328 => x"25732070", 21329 => x"730a0000",
    21330 => x"4d617374", 21331 => x"65722d73", 21332 => x"6c617665",
    21333 => x"2064656c", 21334 => x"61793a20", 21335 => x"20202020",
    21336 => x"20000000", 21337 => x"4d617374", 21338 => x"65722050",
    21339 => x"48592064", 21340 => x"656c6179", 21341 => x"733a2020",
    21342 => x"20202020", 21343 => x"20000000", 21344 => x"54583a20",
    21345 => x"25642070", 21346 => x"732c2052", 21347 => x"583a2025",
    21348 => x"64207073", 21349 => x"0a000000", 21350 => x"536c6176",
    21351 => x"65205048", 21352 => x"59206465", 21353 => x"6c617973",
    21354 => x"3a202020", 21355 => x"20202020", 21356 => x"20000000",
    21357 => x"546f7461", 21358 => x"6c206c69", 21359 => x"6e6b2061",
    21360 => x"73796d6d", 21361 => x"65747279", 21362 => x"3a202020",
    21363 => x"20000000", 21364 => x"25396420", 21365 => x"70730a00",
    21366 => x"4361626c", 21367 => x"65207274", 21368 => x"74206465",
    21369 => x"6c61793a", 21370 => x"20202020", 21371 => x"20202020",
    21372 => x"20000000", 21373 => x"436c6f63", 21374 => x"6b206f66",
    21375 => x"66736574", 21376 => x"3a202020", 21377 => x"20202020",
    21378 => x"20202020", 21379 => x"20000000", 21380 => x"50686173",
    21381 => x"65207365", 21382 => x"74706f69", 21383 => x"6e743a20",
    21384 => x"20202020", 21385 => x"20202020", 21386 => x"20000000",
    21387 => x"536b6577", 21388 => x"3a202020", 21389 => x"20202020",
    21390 => x"20202020", 21391 => x"20202020", 21392 => x"20202020",
    21393 => x"20000000", 21394 => x"55706461", 21395 => x"74652063",
    21396 => x"6f756e74", 21397 => x"65723a20", 21398 => x"20202020",
    21399 => x"20202020", 21400 => x"20000000", 21401 => x"2539640a",
    21402 => x"00000000", 21403 => x"2d2d0000", 21404 => x"756e6b6e",
    21405 => x"6f776e00", 21406 => x"73746174", 21407 => x"73000000",
    21408 => x"1b5b3125", 21409 => x"63000000", 21410 => x"436f6d6d",
    21411 => x"616e6420", 21412 => x"22257322", 21413 => x"3a206572",
    21414 => x"726f7220", 21415 => x"25640a00", 21416 => x"556e7265",
    21417 => x"636f676e", 21418 => x"697a6564", 21419 => x"20636f6d",
    21420 => x"6d616e64", 21421 => x"20222573", 21422 => x"222e0a00",
    21423 => x"77726323", 21424 => x"20000000", 21425 => x"25630000",
    21426 => x"456d7074", 21427 => x"7920696e", 21428 => x"69742073",
    21429 => x"63726970", 21430 => x"742e2e2e", 21431 => x"0a000000",
    21432 => x"65786563", 21433 => x"7574696e", 21434 => x"673a2025",
    21435 => x"730a0000", 21436 => x"57522043", 21437 => x"6f726520",
    21438 => x"6275696c", 21439 => x"643a2025", 21440 => x"7325730a",
    21441 => x"00000000", 21442 => x"2028756e", 21443 => x"73757070",
    21444 => x"6f727465", 21445 => x"64206465", 21446 => x"76656c6f",
    21447 => x"70657220", 21448 => x"6275696c", 21449 => x"64290000",
    21450 => x"4275696c", 21451 => x"743a2025", 21452 => x"73202573",
    21453 => x"20627920", 21454 => x"25730a00", 21455 => x"4275696c",
    21456 => x"7420666f", 21457 => x"72202564", 21458 => x"206b4220",
    21459 => x"52414d2c", 21460 => x"20737461", 21461 => x"636b2069",
    21462 => x"73202564", 21463 => x"20627974", 21464 => x"65730a00",
    21465 => x"5741524e", 21466 => x"494e473a", 21467 => x"20686172",
    21468 => x"64776172", 21469 => x"65207361", 21470 => x"79732025",
    21471 => x"696b4220", 21472 => x"3c3d2052", 21473 => x"414d203c",
    21474 => x"2025696b", 21475 => x"420a0000", 21476 => x"76657200",
    21477 => x"73746172", 21478 => x"74000000", 21479 => x"73746f70",
    21480 => x"00000000", 21481 => x"676d0000", 21482 => x"6d6f6465",
    21483 => x"00000000", 21484 => x"6772616e", 21485 => x"646d6173",
    21486 => x"74657200", 21487 => x"41766169", 21488 => x"6c61626c",
    21489 => x"6520636f", 21490 => x"6d6d616e", 21491 => x"64733a0a",
    21492 => x"00000000", 21493 => x"20202573", 21494 => x"0a000000",
    21495 => x"68656c70", 21496 => x"00000000", 21497 => x"25303278",
    21498 => x"3a253032", 21499 => x"783a2530", 21500 => x"32783a25",
    21501 => x"3032783a", 21502 => x"25303278", 21503 => x"3a253032",
    21504 => x"78000000", 21505 => x"67657400", 21506 => x"67657470",
    21507 => x"00000000", 21508 => x"73657400", 21509 => x"73657470",
    21510 => x"00000000", 21511 => x"4d41432d", 21512 => x"61646472",
    21513 => x"6573733a", 21514 => x"2025730a", 21515 => x"00000000",
    21516 => x"6d616300", 21517 => x"72657365", 21518 => x"74000000",
    21519 => x"20697465", 21520 => x"72617469", 21521 => x"6f6e7320",
    21522 => x"20202020", 21523 => x"7365636f", 21524 => x"6e64732e",
    21525 => x"6d696372", 21526 => x"6f732020", 21527 => x"20206e61",
    21528 => x"6d650a00", 21529 => x"20202539", 21530 => x"6c692020",
    21531 => x"2025396c", 21532 => x"692e2530", 21533 => x"366c6920",
    21534 => x"2025730a", 21535 => x"00000000", 21536 => x"70730000",
    21537 => x"55736167", 21538 => x"653a2072", 21539 => x"65667265",
    21540 => x"7368203c", 21541 => x"7365636f", 21542 => x"6e64733e",
    21543 => x"0a000000", 21544 => x"72656672", 21545 => x"65736800",
    21546 => x"73746174", 21547 => x"69737469", 21548 => x"6373206e",
    21549 => x"6f77206f", 21550 => x"66660a00", 21551 => x"62747300",
    21552 => x"6f666600", 21553 => x"73746174", 21554 => x"00000000",
    21555 => x"57726f6e", 21556 => x"67207061", 21557 => x"72616d65",
    21558 => x"7465720a", 21559 => x"00000000", 21560 => x"65726173",
    21561 => x"65000000", 21562 => x"436f756c", 21563 => x"64206e6f",
    21564 => x"74206572", 21565 => x"61736520", 21566 => x"44420a00",
    21567 => x"61646400", 21568 => x"53465020", 21569 => x"44422069",
    21570 => x"73206675", 21571 => x"6c6c0a00", 21572 => x"49324320",
    21573 => x"6572726f", 21574 => x"720a0000", 21575 => x"53465020",
    21576 => x"64617461", 21577 => x"62617365", 21578 => x"20657272",
    21579 => x"6f722028", 21580 => x"2564290a", 21581 => x"00000000",
    21582 => x"25642053", 21583 => x"46507320", 21584 => x"696e2044",
    21585 => x"420a0000", 21586 => x"73686f77", 21587 => x"00000000",
    21588 => x"53465020", 21589 => x"64617461", 21590 => x"62617365",
    21591 => x"20656d70", 21592 => x"74790a00", 21593 => x"25643a20",
    21594 => x"504e3a00", 21595 => x"20645478", 21596 => x"3a202538",
    21597 => x"64206452", 21598 => x"783a2025", 21599 => x"38642061",
    21600 => x"6c706861", 21601 => x"3a202538", 21602 => x"640a0000",
    21603 => x"6d617463", 21604 => x"68000000", 21605 => x"4e6f2053",
    21606 => x"46502e0a", 21607 => x"00000000", 21608 => x"53465020",
    21609 => x"72656164", 21610 => x"20657272", 21611 => x"6f720a00",
    21612 => x"436f756c", 21613 => x"64206e6f", 21614 => x"74206d61",
    21615 => x"74636820", 21616 => x"746f2044", 21617 => x"420a0000",
    21618 => x"53465020", 21619 => x"6d617463", 21620 => x"6865642c",
    21621 => x"20645478", 21622 => x"3d256420", 21623 => x"6452783d",
    21624 => x"25642061", 21625 => x"6c706861", 21626 => x"3d25640a",
    21627 => x"00000000", 21628 => x"656e6100", 21629 => x"73667000",
    21630 => x"696e6974", 21631 => x"00000000", 21632 => x"636c0000",
    21633 => x"73707300", 21634 => x"67707300", 21635 => x"25642025",
    21636 => x"640a0000", 21637 => x"73646163", 21638 => x"00000000",
    21639 => x"67646163", 21640 => x"00000000", 21641 => x"63686563",
    21642 => x"6b76636f", 21643 => x"00000000", 21644 => x"706c6c00",
    21645 => x"666f7263", 21646 => x"65000000", 21647 => x"466f756e",
    21648 => x"64207068", 21649 => x"61736520", 21650 => x"7472616e",
    21651 => x"73697469", 21652 => x"6f6e2069", 21653 => x"6e204545",
    21654 => x"50524f4d", 21655 => x"3a202564", 21656 => x"70730a00",
    21657 => x"4d656173", 21658 => x"7572696e", 21659 => x"67207432",
    21660 => x"2f743420", 21661 => x"70686173", 21662 => x"65207472",
    21663 => x"616e7369", 21664 => x"74696f6e", 21665 => x"2e2e2e0a",
    21666 => x"00000000", 21667 => x"63616c69", 21668 => x"62726174",
    21669 => x"696f6e00", 21670 => x"73657473", 21671 => x"65630000",
    21672 => x"7365746e", 21673 => x"73656300", 21674 => x"72617700",
    21675 => x"2573202b", 21676 => x"2564206e", 21677 => x"616e6f73",
    21678 => x"65636f6e", 21679 => x"64732e0a", 21680 => x"00000000",
    21681 => x"74696d65", 21682 => x"00000000", 21683 => x"67756900",
    21684 => x"73646200", 21685 => x"4f4e0000", 21686 => x"4f464600",
    21687 => x"656e6162", 21688 => x"6c650000", 21689 => x"64697361",
    21690 => x"626c6500", 21691 => x"70686173", 21692 => x"65207472",
    21693 => x"61636b69", 21694 => x"6e672025", 21695 => x"730a0000",
    21696 => x"70747261", 21697 => x"636b0000", 21698 => x"6c757400",
    21699 => x"6d656173", 21700 => x"00000000", 21701 => x"70636e00",
    21702 => x"25642e25", 21703 => x"642e2564", 21704 => x"2e256400",
    21705 => x"49502d61", 21706 => x"64647265", 21707 => x"73733a20",
    21708 => x"696e2074", 21709 => x"7261696e", 21710 => x"696e670a",
    21711 => x"00000000", 21712 => x"49502d61", 21713 => x"64647265",
    21714 => x"73733a20", 21715 => x"25732028", 21716 => x"66726f6d",
    21717 => x"20626f6f", 21718 => x"7470290a", 21719 => x"00000000",
    21720 => x"49502d61", 21721 => x"64647265", 21722 => x"73733a20",
    21723 => x"25732028", 21724 => x"73746174", 21725 => x"69632061",
    21726 => x"73736967", 21727 => x"6e6d656e", 21728 => x"74290a00",
    21729 => x"69700000", 21730 => x"50505349", 21731 => x"20766572",
    21732 => x"626f7369", 21733 => x"74793a20", 21734 => x"2530386c",
    21735 => x"780a0000", 21736 => x"76657262", 21737 => x"6f736500",
    21738 => x"6465766d", 21739 => x"656d3a20", 21740 => x"7573653a",
    21741 => x"20226465", 21742 => x"766d656d", 21743 => x"203c6164",
    21744 => x"64726573", 21745 => x"733e205b", 21746 => x"3c76616c",
    21747 => x"75653e5d", 21748 => x"220a0000", 21749 => x"25303878",
    21750 => x"203d2025", 21751 => x"3038780a", 21752 => x"00000000",
    21753 => x"64656c61", 21754 => x"79733a20", 21755 => x"7573653a",
    21756 => x"20226465", 21757 => x"6c617973", 21758 => x"205b3c74",
    21759 => x"7864656c", 21760 => x"61793e20", 21761 => x"3c727864",
    21762 => x"656c6179", 21763 => x"3e5d220a", 21764 => x"00000000",
    21765 => x"74783a20", 21766 => x"25692020", 21767 => x"2072783a",
    21768 => x"2025690a", 21769 => x"00000000", 21770 => x"64656c61",
    21771 => x"79730000", 21772 => x"6465766d", 21773 => x"656d0000",
    21774 => x"436f756c", 21775 => x"64206e6f", 21776 => x"74206572",
    21777 => x"61736520", 21778 => x"696e6974", 21779 => x"20736372",
    21780 => x"6970740a", 21781 => x"00000000", 21782 => x"436f756c",
    21783 => x"64206e6f", 21784 => x"74206164", 21785 => x"64207468",
    21786 => x"6520636f", 21787 => x"6d6d616e", 21788 => x"640a0000",
    21789 => x"4f4b2e0a", 21790 => x"00000000", 21791 => x"626f6f74",
    21792 => x"00000000", 21793 => x"25732c20", 21794 => x"25732025",
    21795 => x"642c2025", 21796 => x"642c2025", 21797 => x"3032643a",
    21798 => x"25303264", 21799 => x"3a253032", 21800 => x"64000000",
    21801 => x"25732025", 21802 => x"32642025", 21803 => x"3032643a",
    21804 => x"25303264", 21805 => x"3a253032", 21806 => x"64000000",
    21807 => x"2534642d", 21808 => x"25303264", 21809 => x"2d253032",
    21810 => x"642d2530", 21811 => x"32643a25", 21812 => x"3032643a",
    21813 => x"25303264", 21814 => x"00000000", 21815 => x"1b5b3025",
    21816 => x"643b3325", 21817 => x"646d0000", 21818 => x"1b5b6d00",
    21819 => x"1b5b2564", 21820 => x"3b256466", 21821 => x"00000000",
    21822 => x"1b5b324a", 21823 => x"1b5b313b", 21824 => x"31480000",
    21825 => x"53756e00", 21826 => x"4d6f6e00", 21827 => x"54756500",
    21828 => x"57656400", 21829 => x"54687500", 21830 => x"46726900",
    21831 => x"53617400", 21832 => x"4a616e00", 21833 => x"46656200",
    21834 => x"4d617200", 21835 => x"41707200", 21836 => x"4d617900",
    21837 => x"4a756e00", 21838 => x"4a756c00", 21839 => x"41756700",
    21840 => x"53657000", 21841 => x"4f637400", 21842 => x"4e6f7600",
    21843 => x"44656300", 21844 => x"4c6f6f70", 21845 => x"73207065",
    21846 => x"72206a69", 21847 => x"6666793a", 21848 => x"2025690a",
    21849 => x"00000000", 21850 => x"25733a20", 21851 => x"6e6f2073",
    21852 => x"6f636b65", 21853 => x"7420736c", 21854 => x"6f747320",
    21855 => x"6c656674", 21856 => x"0a000000", 21857 => x"77723000",
    21858 => x"6e65742d", 21859 => x"62680000", 21860 => x"69707634",
    21861 => x"00000000", 21862 => x"61727000", 21863 => x"44697363",
    21864 => x"6f766572", 21865 => x"65642049", 21866 => x"50206164",
    21867 => x"64726573", 21868 => x"73202825", 21869 => x"642e2564",
    21870 => x"2e25642e", 21871 => x"25642921", 21872 => x"0a000000",
    21873 => x"534e4d50", 21874 => x"3a205346", 21875 => x"50207570",
    21876 => x"64617465", 21877 => x"6420696e", 21878 => x"206d656d",
    21879 => x"6f72792c", 21880 => x"20726573", 21881 => x"74617274",
    21882 => x"20505450", 21883 => x"0a000000", 21884 => x"494e5641",
    21885 => x"4c494400", 21886 => x"25642e25", 21887 => x"30346400",
    21888 => x"736e6d70", 21889 => x"00000000", 21890 => x"44656320",
    21891 => x"20362032", 21892 => x"30313620", 21893 => x"31303a30",
    21894 => x"333a3537", 21895 => x"00000000", 21896 => x"30313233",
    21897 => x"34353637", 21898 => x"38396162", 21899 => x"63646566",
    21900 => x"00000000", 21901 => x"49443a20", 21902 => x"25780a00",
    21903 => x"6e6f2070", 21904 => x"66696c74", 21905 => x"65722072",
    21906 => x"756c652d", 21907 => x"73657421", 21908 => x"0a000000",
    21909 => x"7066696c", 21910 => x"7465723a", 21911 => x"2077726f",
    21912 => x"6e67206d", 21913 => x"61676963", 21914 => x"206e756d",
    21915 => x"62657220", 21916 => x"28676f74", 21917 => x"20307825",
    21918 => x"78290a00", 21919 => x"7066696c", 21920 => x"7465723a",
    21921 => x"2077726f", 21922 => x"6e672072", 21923 => x"756c652d",
    21924 => x"7365742c", 21925 => x"2063616e", 21926 => x"27742061",
    21927 => x"70706c79", 21928 => x"0a000000", 21929 => x"696e7661",
    21930 => x"6c696420", 21931 => x"64657363", 21932 => x"72697074",
    21933 => x"6f722040", 21934 => x"2578203d", 21935 => x"2025780a",
    21936 => x"00000000", 21937 => x"5761726e", 21938 => x"696e673a",
    21939 => x"20747820", 21940 => x"6e6f7420", 21941 => x"7465726d",
    21942 => x"696e6174", 21943 => x"65642069", 21944 => x"6e66696e",
    21945 => x"69746520", 21946 => x"6d63723d", 21947 => x"30782578",
    21948 => x"0a000000", 21949 => x"5761726e", 21950 => x"696e673a",
    21951 => x"20747820", 21952 => x"74696d65", 21953 => x"7374616d",
    21954 => x"70206e65", 21955 => x"76657220", 21956 => x"62656361",
    21957 => x"6d652061", 21958 => x"7661696c", 21959 => x"61626c65",
    21960 => x"0a000000", 21961 => x"64657620", 21962 => x"20307825",
    21963 => x"30386c78", 21964 => x"20402025", 21965 => x"30366c78",
    21966 => x"2c202573", 21967 => x"0a000000", 21968 => x"66706761",
    21969 => x"2d617265", 21970 => x"61000000", 21971 => x"4572726f",
    21972 => x"72202564", 21973 => x"20776869", 21974 => x"6c652072",
    21975 => x"65616469", 21976 => x"6e672074", 21977 => x"32347020",
    21978 => x"66726f6d", 21979 => x"2073746f", 21980 => x"72616765",
    21981 => x"0a000000", 21982 => x"74323470", 21983 => x"20726561",
    21984 => x"64206672", 21985 => x"6f6d2073", 21986 => x"746f7261",
    21987 => x"67653a20", 21988 => x"25642070", 21989 => x"730a0000",
    21990 => x"57616974", 21991 => x"696e6720", 21992 => x"666f7220",
    21993 => x"6c696e6b", 21994 => x"2e2e2e0a", 21995 => x"00000000",
    21996 => x"4c6f636b", 21997 => x"696e6720", 21998 => x"504c4c2e",
    21999 => x"2e2e0a00", 22000 => x"43616c69", 22001 => x"62726174",
    22002 => x"696e6720", 22003 => x"52582074", 22004 => x"696d6573",
    22005 => x"74616d70", 22006 => x"65722e2e", 22007 => x"2e0a0000",
    22008 => x"4661696c", 22009 => x"65640000", 22010 => x"53756363",
    22011 => x"65737300", 22012 => x"57726f74", 22013 => x"65206e65",
    22014 => x"77207432", 22015 => x"34702076", 22016 => x"616c7565",
    22017 => x"3a202564", 22018 => x"20707320", 22019 => x"28257329",
    22020 => x"0a000000", 22021 => x"20454e4f", 22022 => x"53504300",
    22023 => x"25732573", 22024 => x"3a000000", 22025 => x"74656d70",
    22026 => x"00000000", 22027 => x"74656d70", 22028 => x"65726174",
    22029 => x"75726500", 22030 => x"55706461", 22031 => x"74652065",
    22032 => x"78697374", 22033 => x"696e6720", 22034 => x"53465020",
    22035 => x"656e7472", 22036 => x"790a0000", 22037 => x"41646469",
    22038 => x"6e67206e", 22039 => x"65772053", 22040 => x"46502065",
    22041 => x"6e747279", 22042 => x"0a000000", 22043 => x"43616e27",
    22044 => x"74207361", 22045 => x"76652070", 22046 => x"65727369",
    22047 => x"7374656e", 22048 => x"74204d41", 22049 => x"43206164",
    22050 => x"64726573", 22051 => x"730a0000", 22052 => x"25733a20",
    22053 => x"5573696e", 22054 => x"67205731", 22055 => x"20736572",
    22056 => x"69616c20", 22057 => x"6e756d62", 22058 => x"65720a00",
    22059 => x"6f666673", 22060 => x"65742025", 22061 => x"34692028",
    22062 => x"30782530", 22063 => x"3378293a", 22064 => x"20253369",
    22065 => x"20283078", 22066 => x"25303278", 22067 => x"290a0000",
    22068 => x"77726974", 22069 => x"65283078", 22070 => x"25782c20",
    22071 => x"2569293a", 22072 => x"20726573", 22073 => x"756c7420",
    22074 => x"3d202569", 22075 => x"0a000000", 22076 => x"72656164",
    22077 => x"28307825", 22078 => x"782c2025", 22079 => x"69293a20",
    22080 => x"72657375", 22081 => x"6c74203d", 22082 => x"2025690a",
    22083 => x"00000000", 22084 => x"64657669", 22085 => x"63652025",
    22086 => x"693a2025", 22087 => x"30387825", 22088 => x"3038780a",
    22089 => x"00000000", 22090 => x"74656d70", 22091 => x"3a202564",
    22092 => x"2e253034", 22093 => x"640a0000", 22094 => x"77310000",
    22095 => x"77317200", 22096 => x"77317700", 22097 => x"3c756e6b",
    22098 => x"6e6f776e", 22099 => x"3e000000", 22100 => x"736f6674",
    22101 => x"706c6c3a", 22102 => x"20697271", 22103 => x"73202564",
    22104 => x"20736571", 22105 => x"20257320", 22106 => x"6d6f6465",
    22107 => x"20256420", 22108 => x"616c6967", 22109 => x"6e6d656e",
    22110 => x"745f7374", 22111 => x"61746520", 22112 => x"25642048",
    22113 => x"4c256420", 22114 => x"4d4c2564", 22115 => x"2048593d",
    22116 => x"2564204d", 22117 => x"593d2564", 22118 => x"2044656c",
    22119 => x"436e743d", 22120 => x"25640a00", 22121 => x"73746172",
    22122 => x"742d6578", 22123 => x"74000000", 22124 => x"77616974",
    22125 => x"2d657874", 22126 => x"00000000", 22127 => x"73746172",
    22128 => x"742d6865", 22129 => x"6c706572", 22130 => x"00000000",
    22131 => x"77616974", 22132 => x"2d68656c", 22133 => x"70657200",
    22134 => x"73746172", 22135 => x"742d6d61", 22136 => x"696e0000",
    22137 => x"77616974", 22138 => x"2d6d6169", 22139 => x"6e000000",
    22140 => x"72656164", 22141 => x"79000000", 22142 => x"636c6561",
    22143 => x"722d6461", 22144 => x"63730000", 22145 => x"77616974",
    22146 => x"2d636c65", 22147 => x"61722d64", 22148 => x"61637300",
    22149 => x"53746163", 22150 => x"6b206f76", 22151 => x"6572666c",
    22152 => x"6f77210a", 22153 => x"00000000", 22154 => x"badc0ffe",
    22155 => x"3b9aca00", 22156 => x"000f4240", 22157 => x"00080030",
    22158 => x"d4a51000", 22159 => x"3b9ac9ff", 22160 => x"c4653600",
    22161 => x"7ffffffe", 22162 => x"80000001", 22163 => x"fff06000",
    22164 => x"0007d000", 22165 => x"41c64e6d", 22166 => x"00010043",
    22167 => x"00010044", 22168 => x"00015180", 22169 => x"83aa7e80",
    22170 => x"7fffffff", 22171 => x"00062000", 22172 => x"005ee000",
    22173 => x"01000001", 22174 => x"11223344", 22175 => x"e0001fff",
    22176 => x"111ee000", 22177 => x"01554000", 22178 => x"0fffffff",
    22179 => x"059682f0", 22180 => x"0ee6b27f", 22181 => x"c0a80001",
    22182 => x"4b002f40", 22183 => x"01312d02", 22184 => x"01312d0a",
    22185 => x"003d0137", 22186 => x"8000001f", 22187 => x"009895b6",
    22188 => x"c4000001", 22189 => x"000186a0", 22190 => x"00ffffff",
    22191 => x"fffdb610", 22192 => x"000249f0", 22193 => x"05f5e100",
    22194 => x"0bebc200", 22195 => x"fa0a1f00", 22196 => x"01312d03",
    22197 => x"5344422d", 22198 => x"011b1900", 22199 => x"00000000",
    22200 => x"70705f64", 22201 => x"6961675f", 22202 => x"70617273",
    22203 => x"65000000", 22204 => x"00000000", 22205 => x"00013878",
    22206 => x"00013884", 22207 => x"00013894", 22208 => x"000138a0",
    22209 => x"000138ac", 22210 => x"000138b8", 22211 => x"000138c4",
    22212 => x"000014dc", 22213 => x"0000154c", 22214 => x"00001804",
    22215 => x"00001804", 22216 => x"00001804", 22217 => x"00001804",
    22218 => x"00001804", 22219 => x"00001804", 22220 => x"000015c8",
    22221 => x"00001638", 22222 => x"00001804", 22223 => x"000016cc",
    22224 => x"000017d8", 22225 => x"77727063", 22226 => x"5f74696d",
    22227 => x"655f6164", 22228 => x"6a757374", 22229 => x"5f6f6666",
    22230 => x"73657400", 22231 => x"77725f73", 22232 => x"31000000",
    22233 => x"77727063", 22234 => x"5f74696d", 22235 => x"655f6164",
    22236 => x"6a757374", 22237 => x"00000000", 22238 => x"77727063",
    22239 => x"5f74696d", 22240 => x"655f7365", 22241 => x"74000000",
    22242 => x"77727063", 22243 => x"5f74696d", 22244 => x"655f6765",
    22245 => x"74000000", 22246 => x"77727063", 22247 => x"5f6e6574",
    22248 => x"5f73656e", 22249 => x"64000000", 22250 => x"77725f75",
    22251 => x"6e706163", 22252 => x"6b5f616e", 22253 => x"6e6f756e",
    22254 => x"63650000", 22255 => x"77725f70", 22256 => x"61636b5f",
    22257 => x"616e6e6f", 22258 => x"756e6365", 22259 => x"00000000",
    22260 => x"77725f68", 22261 => x"616e646c", 22262 => x"655f666f",
    22263 => x"6c6c6f77", 22264 => x"75700000", 22265 => x"77725f68",
    22266 => x"616e646c", 22267 => x"655f616e", 22268 => x"6e6f756e",
    22269 => x"63650000", 22270 => x"77725f65", 22271 => x"78656375",
    22272 => x"74655f73", 22273 => x"6c617665", 22274 => x"00000000",
    22275 => x"77725f68", 22276 => x"616e646c", 22277 => x"655f7265",
    22278 => x"73700000", 22279 => x"77725f6e", 22280 => x"65775f73",
    22281 => x"6c617665", 22282 => x"00000000", 22283 => x"77725f6d",
    22284 => x"61737465", 22285 => x"725f6d73", 22286 => x"67000000",
    22287 => x"77725f6c", 22288 => x"69737465", 22289 => x"6e696e67",
    22290 => x"00000000", 22291 => x"77725f6f", 22292 => x"70656e00",
    22293 => x"77725f69", 22294 => x"6e697400", 22295 => x"00002ddc",
    22296 => x"00002e04", 22297 => x"00002e24", 22298 => x"00002e94",
    22299 => x"00002eb4", 22300 => x"00002ed0", 22301 => x"00002ef0",
    22302 => x"00002f7c", 22303 => x"00002f9c", 22304 => x"77725f63",
    22305 => x"616c6962", 22306 => x"72617469", 22307 => x"6f6e0000",
    22308 => x"00004420", 22309 => x"00004408", 22310 => x"00004448",
    22311 => x"00004554", 22312 => x"0000449c", 22313 => x"000141e0",
    22314 => x"00014314", 22315 => x"00014320", 22316 => x"0001432c",
    22317 => x"00014338", 22318 => x"00014344", 22319 => x"77725f73",
    22320 => x"6572766f", 22321 => x"5f757064", 22322 => x"61746500",
    22323 => x"70705f69", 22324 => x"6e697469", 22325 => x"616c697a",
    22326 => x"696e6700", 22327 => x"73745f63", 22328 => x"6f6d5f73",
    22329 => x"6c617665", 22330 => x"5f68616e", 22331 => x"646c655f",
    22332 => x"666f6c6c", 22333 => x"6f777570", 22334 => x"00000000",
    22335 => x"626d635f", 22336 => x"64617461", 22337 => x"7365745f",
    22338 => x"636d7000", 22339 => x"626d635f", 22340 => x"73746174",
    22341 => x"655f6465", 22342 => x"63697369", 22343 => x"6f6e0000",
    22344 => x"63466965", 22345 => x"6c645f74", 22346 => x"6f5f5469",
    22347 => x"6d65496e", 22348 => x"7465726e", 22349 => x"616c0000",
    22350 => x"00014e70", 22351 => x"00014fb0", 22352 => x"0001435c",
    22353 => x"00013e74", 22354 => x"0000001f", 22355 => x"0000001c",
    22356 => x"0000001f", 22357 => x"0000001e", 22358 => x"0000001f",
    22359 => x"0000001e", 22360 => x"0000001f", 22361 => x"0000001f",
    22362 => x"0000001e", 22363 => x"0000001f", 22364 => x"0000001e",
    22365 => x"0000001f", 22366 => x"0000001f", 22367 => x"0000001d",
    22368 => x"0000001f", 22369 => x"0000001e", 22370 => x"0000001f",
    22371 => x"0000001e", 22372 => x"0000001f", 22373 => x"0000001f",
    22374 => x"0000001e", 22375 => x"0000001f", 22376 => x"0000001e",
    22377 => x"0000001f", 22378 => x"00015504", 22379 => x"00015508",
    22380 => x"0001550c", 22381 => x"00015510", 22382 => x"00015514",
    22383 => x"00015518", 22384 => x"0001551c", 22385 => x"00015520",
    22386 => x"00015524", 22387 => x"00015528", 22388 => x"0001552c",
    22389 => x"00015530", 22390 => x"00015534", 22391 => x"00015538",
    22392 => x"0001553c", 22393 => x"00015540", 22394 => x"00015544",
    22395 => x"00015548", 22396 => x"0001554c", 22397 => x"70747064",
    22398 => x"5f6e6574", 22399 => x"69665f63", 22400 => x"72656174",
    22401 => x"655f736f", 22402 => x"636b6574", 22403 => x"00000000",
    22404 => x"0000b7d4", 22405 => x"0000b7e4", 22406 => x"0000b848",
    22407 => x"0000b848", 22408 => x"0000b7f4", 22409 => x"0000b848",
    22410 => x"0000b848", 22411 => x"30ff0201", 22412 => x"fa040670",
    22413 => x"75626c69", 22414 => x"63fdff02", 22415 => x"f90201fc",
    22416 => x"0201fb30", 22417 => x"ff30ff06", 22418 => x"6765745f",
    22419 => x"70657273", 22420 => x"69737465", 22421 => x"6e745f6d",
    22422 => x"61630000", 22423 => x"000000c8", 22424 => x"000039d0",
    22425 => x"00010d78", 22426 => x"00010dfc", 22427 => x"00010e34",
    22428 => x"00010eb4", 22429 => x"00010f40", 22430 => x"00010f58",
    22431 => x"00010e58", 22432 => x"00010da0", 22433 => x"00010cfc",
    22434 => x"00010d30", 22435 => x"00000000", 22436 => x"00000000",
    22437 => x"00000000", 22438 => x"00000000", 22439 => x"00000001",
    22440 => x"00000001", 22441 => x"00000001", 22442 => x"00000001",
    22443 => x"00000000", 22444 => x"00000000", 22445 => x"00000000",
    22446 => x"0000ece8", 22447 => x"0000ece8", 22448 => x"00000000",
    22449 => x"0000d9d0", 22450 => x"00000000", 22451 => x"00011abc",
    22452 => x"00011adc", 22453 => x"00011ae8", 22454 => x"00011af8",
    22455 => x"00011b18", 22456 => x"00011b28", 22457 => x"00011b7c",
    22458 => x"00011b40", 22459 => x"00011a50", 22460 => x"00011a94",
    22461 => x"00000001", 22462 => x"000159a4", 22463 => x"00000002",
    22464 => x"000159b0", 22465 => x"00000003", 22466 => x"000159bc",
    22467 => x"00000004", 22468 => x"000159cc", 22469 => x"00000005",
    22470 => x"000159d8", 22471 => x"00000006", 22472 => x"000159e4",
    22473 => x"00000007", 22474 => x"00013e4c", 22475 => x"00000008",
    22476 => x"000159f0", 22477 => x"00000009", 22478 => x"000159f8",
    22479 => x"0000000a", 22480 => x"00015a04", 22481 => x"00000000",
    22482 => x"00000000", 22483 => x"00000000", 22484 => x"00000000",
    22485 => x"00000000", 22486 => x"00000000", 22487 => x"00010000",
    22488 => x"00000000", 22489 => x"00000000", 22490 => x"00000000",
    22491 => x"00020100", 22492 => x"00000000", 22493 => x"00000000",
    22494 => x"00000000", 22495 => x"00030101", 22496 => x"00000000",
    22497 => x"00000000", 22498 => x"00000000", 22499 => x"00040201",
    22500 => x"01000000", 22501 => x"00000000", 22502 => x"00000000",
    22503 => x"00050201", 22504 => x"01010000", 22505 => x"00000000",
    22506 => x"00000000", 22507 => x"00060302", 22508 => x"01010100",
    22509 => x"00000000", 22510 => x"00000000", 22511 => x"00070302",
    22512 => x"01010101", 22513 => x"00000000", 22514 => x"00000000",
    22515 => x"00080402", 22516 => x"02010101", 22517 => x"01000000",
    22518 => x"00000000", 22519 => x"00090403", 22520 => x"02010101",
    22521 => x"01010000", 22522 => x"00000000", 22523 => x"000a0503",
    22524 => x"02020101", 22525 => x"01010100", 22526 => x"00000000",
    22527 => x"000b0503", 22528 => x"02020101", 22529 => x"01010101",
    22530 => x"00000000", 22531 => x"000c0604", 22532 => x"03020201",
    22533 => x"01010101", 22534 => x"01000000", 22535 => x"000d0604",
    22536 => x"03020201", 22537 => x"01010101", 22538 => x"01010000",
    22539 => x"000e0704", 22540 => x"03020202", 22541 => x"01010101",
    22542 => x"01010100", 22543 => x"000f0705", 22544 => x"03030202",
    22545 => x"01010101", 22546 => x"01010101", 22547 => x"fefefeff",
    22548 => x"80808080", 22549 => x"00202020", 22550 => x"20202020",
    22551 => x"20202828", 22552 => x"28282820", 22553 => x"20202020",
    22554 => x"20202020", 22555 => x"20202020", 22556 => x"20202020",
    22557 => x"20881010", 22558 => x"10101010", 22559 => x"10101010",
    22560 => x"10101010", 22561 => x"10040404", 22562 => x"04040404",
    22563 => x"04040410", 22564 => x"10101010", 22565 => x"10104141",
    22566 => x"41414141", 22567 => x"01010101", 22568 => x"01010101",
    22569 => x"01010101", 22570 => x"01010101", 22571 => x"01010101",
    22572 => x"10101010", 22573 => x"10104242", 22574 => x"42424242",
    22575 => x"02020202", 22576 => x"02020202", 22577 => x"02020202",
    22578 => x"02020202", 22579 => x"02020202", 22580 => x"10101010",
    22581 => x"20000000", 22582 => x"00000000", 22583 => x"00000000",
    22584 => x"00000000", 22585 => x"00000000", 22586 => x"00000000",
    22587 => x"00000000", 22588 => x"00000000", 22589 => x"00000000",
    22590 => x"00000000", 22591 => x"00000000", 22592 => x"00000000",
    22593 => x"00000000", 22594 => x"00000000", 22595 => x"00000000",
    22596 => x"00000000", 22597 => x"00000000", 22598 => x"00000000",
    22599 => x"00000000", 22600 => x"00000000", 22601 => x"00000000",
    22602 => x"00000000", 22603 => x"00000000", 22604 => x"00000000",
    22605 => x"00000000", 22606 => x"00000000", 22607 => x"00000000",
    22608 => x"00000000", 22609 => x"00000000", 22610 => x"00000000",
    22611 => x"00000000", 22612 => x"00000000", 22613 => x"00000000",
    22614 => x"000172f0", 22615 => x"00017310", 22616 => x"00017320",
    22617 => x"00017330", 22618 => x"000003e8", 22619 => x"00000001",
    22620 => x"00000955", 22621 => x"ffffffff", 22622 => x"00000000",
    22623 => x"00000000", 22624 => x"00000000", 22625 => x"00000000",
    22626 => x"00000000", 22627 => x"00000000", 22628 => x"00000000",
    22629 => x"00000000", 22630 => x"000164ec", 22631 => x"0001660c",
    22632 => x"000165f0", 22633 => x"000175a0", 22634 => x"00017620",
    22635 => x"00000000", 22636 => x"00000000", 22637 => x"00000000",
    22638 => x"00000000", 22639 => x"00000000", 22640 => x"00000000",
    22641 => x"00000000", 22642 => x"00000000", 22643 => x"00000000",
    22644 => x"00000000", 22645 => x"00000000", 22646 => x"00000000",
    22647 => x"00000000", 22648 => x"00000000", 22649 => x"00000000",
    22650 => x"00000000", 22651 => x"00000000", 22652 => x"00000000",
    22653 => x"00000000", 22654 => x"00000000", 22655 => x"00000000",
    22656 => x"00000000", 22657 => x"00000000", 22658 => x"00000000",
    22659 => x"00000000", 22660 => x"00000000", 22661 => x"00000000",
    22662 => x"00000000", 22663 => x"00000000", 22664 => x"00000000",
    22665 => x"00000000", 22666 => x"00000000", 22667 => x"00000000",
    22668 => x"00000000", 22669 => x"00000000", 22670 => x"00000000",
    22671 => x"00000000", 22672 => x"00000000", 22673 => x"00000000",
    22674 => x"00000000", 22675 => x"00000000", 22676 => x"00000000",
    22677 => x"00000000", 22678 => x"00000000", 22679 => x"00000000",
    22680 => x"00000000", 22681 => x"00000000", 22682 => x"00000000",
    22683 => x"00000000", 22684 => x"00000000", 22685 => x"00000000",
    22686 => x"00000000", 22687 => x"00000000", 22688 => x"00000000",
    22689 => x"00000000", 22690 => x"00000000", 22691 => x"00000000",
    22692 => x"00000000", 22693 => x"00000000", 22694 => x"00000000",
    22695 => x"00000000", 22696 => x"00000000", 22697 => x"00000000",
    22698 => x"00000000", 22699 => x"00000000", 22700 => x"00000000",
    22701 => x"00000000", 22702 => x"00000000", 22703 => x"00000000",
    22704 => x"00000000", 22705 => x"00000000", 22706 => x"00000000",
    22707 => x"00000000", 22708 => x"00000000", 22709 => x"00000000",
    22710 => x"00000000", 22711 => x"00000000", 22712 => x"00000000",
    22713 => x"00000000", 22714 => x"00000000", 22715 => x"00000000",
    22716 => x"00000000", 22717 => x"00000000", 22718 => x"00000000",
    22719 => x"00000000", 22720 => x"00000000", 22721 => x"00000000",
    22722 => x"00000000", 22723 => x"00000000", 22724 => x"00000000",
    22725 => x"00000000", 22726 => x"00000000", 22727 => x"00000000",
    22728 => x"00000000", 22729 => x"00000000", 22730 => x"00000000",
    22731 => x"00000000", 22732 => x"00000000", 22733 => x"00000000",
    22734 => x"00000000", 22735 => x"00000000", 22736 => x"00000000",
    22737 => x"00000000", 22738 => x"00000000", 22739 => x"00000000",
    22740 => x"00000000", 22741 => x"00000000", 22742 => x"00000000",
    22743 => x"00000000", 22744 => x"00000000", 22745 => x"00000000",
    22746 => x"00000000", 22747 => x"00000000", 22748 => x"00000000",
    22749 => x"00000000", 22750 => x"00000000", 22751 => x"00000000",
    22752 => x"00000000", 22753 => x"00000000", 22754 => x"00000000",
    22755 => x"00000000", 22756 => x"00000000", 22757 => x"00000000",
    22758 => x"00000000", 22759 => x"00000000", 22760 => x"00000000",
    22761 => x"00000000", 22762 => x"00000000", 22763 => x"00000000",
    22764 => x"00000000", 22765 => x"00000000", 22766 => x"00000000",
    22767 => x"00000000", 22768 => x"00000000", 22769 => x"00000000",
    22770 => x"00000000", 22771 => x"00000000", 22772 => x"00000000",
    22773 => x"00000000", 22774 => x"00000000", 22775 => x"00000000",
    22776 => x"00000000", 22777 => x"00000000", 22778 => x"00000000",
    22779 => x"00000000", 22780 => x"00000000", 22781 => x"00000000",
    22782 => x"00000000", 22783 => x"00000000", 22784 => x"00000000",
    22785 => x"00000000", 22786 => x"00000000", 22787 => x"00000000",
    22788 => x"00000000", 22789 => x"00000000", 22790 => x"00000000",
    22791 => x"00000000", 22792 => x"00000000", 22793 => x"00000000",
    22794 => x"00000000", 22795 => x"00000000", 22796 => x"00000000",
    22797 => x"00000000", 22798 => x"00000000", 22799 => x"00000000",
    22800 => x"00016534", 22801 => x"00000000", 22802 => x"00000000",
    22803 => x"00000000", 22804 => x"00000000", 22805 => x"00000000",
    22806 => x"00000000", 22807 => x"00000000", 22808 => x"00000000",
    22809 => x"00000000", 22810 => x"00000000", 22811 => x"00000000",
    22812 => x"00000000", 22813 => x"00000000", 22814 => x"00000000",
    22815 => x"00000000", 22816 => x"00000000", 22817 => x"00000000",
    22818 => x"00000000", 22819 => x"00000000", 22820 => x"00000000",
    22821 => x"00000000", 22822 => x"00000000", 22823 => x"00000000",
    22824 => x"00000000", 22825 => x"00000000", 22826 => x"00013954",
    22827 => x"00013954", 22828 => x"00000000", 22829 => x"00000001",
    22830 => x"00000000", 22831 => x"00000000", 22832 => x"00000000",
    22833 => x"00000000", 22834 => x"00000000", 22835 => x"00000000",
    22836 => x"00000000", 22837 => x"00000000", 22838 => x"00000000",
    22839 => x"00000000", 22840 => x"00000000", 22841 => x"00000000",
    22842 => x"00000000", 22843 => x"00016178", 22844 => x"000176a0",
    22845 => x"00000000", 22846 => x"000176e0", 22847 => x"000176fc",
    22848 => x"0001772c", 22849 => x"0001774c", 22850 => x"00000000",
    22851 => x"00000000", 22852 => x"00000000", 22853 => x"00000000",
    22854 => x"00000000", 22855 => x"00000000", 22856 => x"00000000",
    22857 => x"00000000", 22858 => x"00000000", 22859 => x"00017770",
    22860 => x"000003e8", 22861 => x"00000000", 22862 => x"00000000",
    22863 => x"00000000", 22864 => x"00000000", 22865 => x"00016548",
    22866 => x"000165b4", 22867 => x"00000000", 22868 => x"00000000",
    22869 => x"00000000", 22870 => x"00000000", 22871 => x"00000000",
    22872 => x"00000000", 22873 => x"00000000", 22874 => x"00000000",
    22875 => x"00000000", 22876 => x"00000000", 22877 => x"00000000",
    22878 => x"00000000", 22879 => x"00000000", 22880 => x"00000000",
    22881 => x"00000000", 22882 => x"00000000", 22883 => x"00000000",
    22884 => x"00000000", 22885 => x"00000000", 22886 => x"00000000",
    22887 => x"00000000", 22888 => x"00000000", 22889 => x"00000000",
    22890 => x"00000000", 22891 => x"00000000", 22892 => x"00000000",
    22893 => x"00000a58", 22894 => x"00000a8c", 22895 => x"00000b0c",
    22896 => x"00000b14", 22897 => x"00000b6c", 22898 => x"00000b98",
    22899 => x"00000bf0", 22900 => x"00000c14", 22901 => x"00000cd8",
    22902 => x"00000ce0", 22903 => x"00000ce8", 22904 => x"00000d4c",
    22905 => x"00000d68", 22906 => x"00000b38", 22907 => x"00000000",
    22908 => x"00001c8c", 22909 => x"00001c10", 22910 => x"00001bb4",
    22911 => x"00001b5c", 22912 => x"00000000", 22913 => x"00000000",
    22914 => x"00001b2c", 22915 => x"00001f18", 22916 => x"00001ef8",
    22917 => x"00001e28", 22918 => x"00001d0c", 22919 => x"00000000",
    22920 => x"00000000", 22921 => x"00000000", 22922 => x"00000000",
    22923 => x"00000000", 22924 => x"00000000", 22925 => x"00000000",
    22926 => x"00000000", 22927 => x"00000000", 22928 => x"00000000",
    22929 => x"00000000", 22930 => x"00000200", 22931 => x"00000000",
    22932 => x"00017880", 22933 => x"00000001", 22934 => x"00013e34",
    22935 => x"00004748", 22936 => x"00000002", 22937 => x"00013e44",
    22938 => x"00004914", 22939 => x"00000003", 22940 => x"00013e4c",
    22941 => x"000049d0", 22942 => x"00000004", 22943 => x"00013e58",
    22944 => x"000049e0", 22945 => x"00000006", 22946 => x"0001435c",
    22947 => x"00004b8c", 22948 => x"00000008", 22949 => x"00013e64",
    22950 => x"00004ecc", 22951 => x"00000009", 22952 => x"00013e74",
    22953 => x"00004f40", 22954 => x"00000064", 22955 => x"00013e7c",
    22956 => x"00002814", 22957 => x"00000066", 22958 => x"00013e94",
    22959 => x"0000298c", 22960 => x"00000065", 22961 => x"00013ea8",
    22962 => x"00002ab8", 22963 => x"00000067", 22964 => x"00013ec0",
    22965 => x"00002bbc", 22966 => x"00000068", 22967 => x"00013ed8",
    22968 => x"00002ce8", 22969 => x"00000069", 22970 => x"00013ee8",
    22971 => x"00003004", 22972 => x"0000006a", 22973 => x"00013ef8",
    22974 => x"00003118", 22975 => x"0000006b", 22976 => x"00013f0c",
    22977 => x"0000329c", 22978 => x"00000000", 22979 => x"00000000",
    22980 => x"00000000", 22981 => x"00000001", 22982 => x"00013e34",
    22983 => x"00004748", 22984 => x"00000002", 22985 => x"00013e44",
    22986 => x"00004914", 22987 => x"00000003", 22988 => x"00013e4c",
    22989 => x"000049d0", 22990 => x"00000004", 22991 => x"00013e58",
    22992 => x"000049e0", 22993 => x"00000005", 22994 => x"00014358",
    22995 => x"00004af8", 22996 => x"00000006", 22997 => x"0001435c",
    22998 => x"00004b8c", 22999 => x"00000007", 23000 => x"00014364",
    23001 => x"00004e08", 23002 => x"00000008", 23003 => x"00013e64",
    23004 => x"00004ecc", 23005 => x"00000009", 23006 => x"00013e74",
    23007 => x"00004f40", 23008 => x"00000000", 23009 => x"00000000",
    23010 => x"00000000", 23011 => x"00002218", 23012 => x"00002138",
    23013 => x"00000000", 23014 => x"000020f0", 23015 => x"000025b0",
    23016 => x"00002568", 23017 => x"0000247c", 23018 => x"00002060",
    23019 => x"00001fd4", 23020 => x"00002404", 23021 => x"0000238c",
    23022 => x"00002324", 23023 => x"000022b8", 23024 => x"00000001",
    23025 => x"00014570", 23026 => x"00014578", 23027 => x"00014584",
    23028 => x"00014590", 23029 => x"00000000", 23030 => x"00000000",
    23031 => x"00000000", 23032 => x"00000000", 23033 => x"000145b4",
    23034 => x"0001459c", 23035 => x"000145a8", 23036 => x"000145c0",
    23037 => x"000145cc", 23038 => x"000145d8", 23039 => x"00000000",
    23040 => x"00000000", 23041 => x"00014900", 23042 => x"00014910",
    23043 => x"0001491c", 23044 => x"00014930", 23045 => x"00014944",
    23046 => x"00014954", 23047 => x"00014960", 23048 => x"0001496c",
    23049 => x"bbfef060", 23050 => x"00000000", 23051 => x"00000000",
    23052 => x"00000000", 23053 => x"00000000", 23054 => x"00000000",
    23055 => x"00000000", 23056 => x"00000000", 23057 => x"00000000",
    23058 => x"00000000", 23059 => x"00000000", 23060 => x"00000000",
    23061 => x"00000000", 23062 => x"00000001", 23063 => x"00000000",
    23064 => x"000a03e8", 23065 => x"00060100", 23066 => x"80800000",
    23067 => x"00000000", 23068 => x"00016178", 23069 => x"00000000",
    23070 => x"00000000", 23071 => x"00000000", 23072 => x"00000000",
    23073 => x"00000000", 23074 => x"00000000", 23075 => x"00000000",
    23076 => x"00000000", 23077 => x"00000000", 23078 => x"00000000",
    23079 => x"00000200", 23080 => x"00000000", 23081 => x"00017dac",
    23082 => x"00000000", 23083 => x"00000000", 23084 => x"00000000",
    23085 => x"00000000", 23086 => x"00000000", 23087 => x"00000000",
    23088 => x"00000000", 23089 => x"00000000", 23090 => x"00000000",
    23091 => x"00000000", 23092 => x"00000060", 23093 => x"00000000",
    23094 => x"00017fac", 23095 => x"00000000", 23096 => x"00000000",
    23097 => x"00000000", 23098 => x"00000000", 23099 => x"00000000",
    23100 => x"00000000", 23101 => x"00000000", 23102 => x"00000000",
    23103 => x"00000000", 23104 => x"00000000", 23105 => x"00000080",
    23106 => x"00000000", 23107 => x"0001800c", 23108 => x"00000000",
    23109 => x"00000000", 23110 => x"00000000", 23111 => x"00000000",
    23112 => x"00000000", 23113 => x"00000000", 23114 => x"00000000",
    23115 => x"00000000", 23116 => x"00000000", 23117 => x"00000000",
    23118 => x"00000080", 23119 => x"00000000", 23120 => x"00018090",
    23121 => x"63757465", 23122 => x"70636e00", 23123 => x"00000000",
    23124 => x"00000000", 23125 => x"00000000", 23126 => x"00000000",
    23127 => x"00000000", 23128 => x"00000000", 23129 => x"00016a28",
    23130 => x"0000bd24", 23131 => x"00016a34", 23132 => x"09000000",
    23133 => x"00016a98", 23134 => x"0000bd24", 23135 => x"00016aa4",
    23136 => x"09000000", 23137 => x"00016af4", 23138 => x"0000bb14",
    23139 => x"00016b00", 23140 => x"0a000000", 23141 => x"00016b3c",
    23142 => x"0000bd24", 23143 => x"00016b48", 23144 => x"09000000",
    23145 => x"00016c10", 23146 => x"0000bd24", 23147 => x"00016c1c",
    23148 => x"09000000", 23149 => x"00016d84", 23150 => x"0000bd24",
    23151 => x"00016d90", 23152 => x"09000000", 23153 => x"00016e1c",
    23154 => x"0000bd24", 23155 => x"00016e28", 23156 => x"09000000",
    23157 => x"00016ea0", 23158 => x"0000bb14", 23159 => x"00016eac",
    23160 => x"0a000000", 23161 => x"00000000", 23162 => x"00000000",
    23163 => x"00000000", 23164 => x"00000000", 23165 => x"00000000",
    23166 => x"00000000", 23167 => x"00000000", 23168 => x"00000000",
    23169 => x"00000000", 23170 => x"00000000", 23171 => x"00000000",
    23172 => x"00000000", 23173 => x"00000000", 23174 => x"00000000",
    23175 => x"00000100", 23176 => x"00000000", 23177 => x"00018138",
    23178 => x"2b060104", 23179 => x"01606501", 23180 => x"01000000",
    23181 => x"00016f10", 23182 => x"0000c2a0", 23183 => x"00000000",
    23184 => x"00016944", 23185 => x"02040020", 23186 => x"00016f14",
    23187 => x"0000c274", 23188 => x"00000000", 23189 => x"00016158",
    23190 => x"02040004", 23191 => x"00016f18", 23192 => x"0000c274",
    23193 => x"00000000", 23194 => x"00016164", 23195 => x"02040004",
    23196 => x"00016f1c", 23197 => x"0000c274", 23198 => x"00000000",
    23199 => x"00016f20", 23200 => x"02040004", 23201 => x"00000000",
    23202 => x"00000000", 23203 => x"00000000", 23204 => x"00000000",
    23205 => x"00000000", 23206 => x"2b060104", 23207 => x"01606501",
    23208 => x"02000000", 23209 => x"00016f24", 23210 => x"0000c638",
    23211 => x"00000000", 23212 => x"00000004", 23213 => x"02460001",
    23214 => x"00016f28", 23215 => x"0000c638", 23216 => x"00000000",
    23217 => x"00000005", 23218 => x"02040001", 23219 => x"00016f2c",
    23220 => x"0000c638", 23221 => x"00000000", 23222 => x"00000002",
    23223 => x"02430001", 23224 => x"00000000", 23225 => x"00000000",
    23226 => x"00000000", 23227 => x"00000000", 23228 => x"00000000",
    23229 => x"2b060104", 23230 => x"01606501", 23231 => x"03010000",
    23232 => x"00016f30", 23233 => x"0000c508", 23234 => x"00000000",
    23235 => x"00000000", 23236 => x"01040001", 23237 => x"00016f34",
    23238 => x"0000c508", 23239 => x"00000000", 23240 => x"00000000",
    23241 => x"01040001", 23242 => x"00000000", 23243 => x"00000000",
    23244 => x"00000000", 23245 => x"00000000", 23246 => x"00000000",
    23247 => x"2b060104", 23248 => x"01606501", 23249 => x"04000000",
    23250 => x"00016f38", 23251 => x"0000c2a0", 23252 => x"00000000",
    23253 => x"000172c8", 23254 => x"02020004", 23255 => x"00016f3c",
    23256 => x"0000c2a0", 23257 => x"00000000", 23258 => x"000172cc",
    23259 => x"02410004", 23260 => x"00016f40", 23261 => x"0000c2a0",
    23262 => x"00000000", 23263 => x"000172d0", 23264 => x"02020004",
    23265 => x"00016f44", 23266 => x"0000c2a0", 23267 => x"00000000",
    23268 => x"000172d4", 23269 => x"02020004", 23270 => x"00016f48",
    23271 => x"0000c2a0", 23272 => x"00000000", 23273 => x"000172d8",
    23274 => x"02410004", 23275 => x"00016f4c", 23276 => x"0000c2a0",
    23277 => x"00000000", 23278 => x"000172dc", 23279 => x"02410004",
    23280 => x"00016f50", 23281 => x"0000c2a0", 23282 => x"00000000",
    23283 => x"000172e0", 23284 => x"02020004", 23285 => x"00016f54",
    23286 => x"0000c2a0", 23287 => x"00000000", 23288 => x"000172e4",
    23289 => x"02020004", 23290 => x"00016f58", 23291 => x"0000c2a0",
    23292 => x"00000000", 23293 => x"000172e8", 23294 => x"02410004",
    23295 => x"00000000", 23296 => x"00000000", 23297 => x"00000000",
    23298 => x"00000000", 23299 => x"00000000", 23300 => x"2b060104",
    23301 => x"01606501", 23302 => x"05000000", 23303 => x"00016f5c",
    23304 => x"0000c274", 23305 => x"00000000", 23306 => x"00018114",
    23307 => x"02021404", 23308 => x"00016f60", 23309 => x"0000c1e8",
    23310 => x"00000000", 23311 => x"00018114", 23312 => x"0202e808",
    23313 => x"00016f64", 23314 => x"0000c1e8", 23315 => x"00000000",
    23316 => x"00018114", 23317 => x"0202e008", 23318 => x"00016f68",
    23319 => x"0000c274", 23320 => x"00000000", 23321 => x"00018114",
    23322 => x"0246a008", 23323 => x"00016f6c", 23324 => x"0000c274",
    23325 => x"00000000", 23326 => x"00018114", 23327 => x"0241b804",
    23328 => x"00016f70", 23329 => x"0000c0e8", 23330 => x"00000000",
    23331 => x"00000001", 23332 => x"02460001", 23333 => x"00016f74",
    23334 => x"0000c274", 23335 => x"00000000", 23336 => x"00018114",
    23337 => x"02021804", 23338 => x"00016f78", 23339 => x"0000c274",
    23340 => x"00000000", 23341 => x"00018114", 23342 => x"02021c04",
    23343 => x"00016f7c", 23344 => x"0000c274", 23345 => x"00000000",
    23346 => x"00018114", 23347 => x"02022004", 23348 => x"00016f80",
    23349 => x"0000c274", 23350 => x"00000000", 23351 => x"00018114",
    23352 => x"02022404", 23353 => x"00016f84", 23354 => x"0000c274",
    23355 => x"00000000", 23356 => x"00018114", 23357 => x"0241f004",
    23358 => x"00016f88", 23359 => x"0000c274", 23360 => x"00000000",
    23361 => x"00018114", 23362 => x"0241f404", 23363 => x"00016f8c",
    23364 => x"0000c274", 23365 => x"00000000", 23366 => x"00018114",
    23367 => x"0241f804", 23368 => x"00016f90", 23369 => x"0000c0e8",
    23370 => x"00000000", 23371 => x"00000002", 23372 => x"02460001",
    23373 => x"00016f94", 23374 => x"0000c2a0", 23375 => x"00000000",
    23376 => x"000164e4", 23377 => x"02410004", 23378 => x"00016f98",
    23379 => x"0000c2a0", 23380 => x"00000000", 23381 => x"000164e8",
    23382 => x"02410004", 23383 => x"00016f9c", 23384 => x"0000c274",
    23385 => x"00000000", 23386 => x"00018114", 23387 => x"02022804",
    23388 => x"00000000", 23389 => x"00000000", 23390 => x"00000000",
    23391 => x"00000000", 23392 => x"00000000", 23393 => x"2b060104",
    23394 => x"01606501", 23395 => x"06000000", 23396 => x"00016fa0",
    23397 => x"0000c2a0", 23398 => x"0000c328", 23399 => x"00018238",
    23400 => x"02020004", 23401 => x"00016fa4", 23402 => x"0000c2a0",
    23403 => x"0000c388", 23404 => x"0001823c", 23405 => x"02020004",
    23406 => x"00016fa8", 23407 => x"0000c2a0", 23408 => x"0000baf0",
    23409 => x"00018118", 23410 => x"02040010", 23411 => x"00016fac",
    23412 => x"0000c2a0", 23413 => x"0000baf0", 23414 => x"0001812c",
    23415 => x"02020004", 23416 => x"00016fb0", 23417 => x"0000c2a0",
    23418 => x"0000baf0", 23419 => x"00018130", 23420 => x"02020004",
    23421 => x"00016fb4", 23422 => x"0000c2a0", 23423 => x"0000baf0",
    23424 => x"00018128", 23425 => x"02020004", 23426 => x"00000000",
    23427 => x"00000000", 23428 => x"00000000", 23429 => x"00000000",
    23430 => x"00000000", 23431 => x"2b060104", 23432 => x"01606501",
    23433 => x"07000000", 23434 => x"00016fb8", 23435 => x"0000c2c8",
    23436 => x"00000000", 23437 => x"00000001", 23438 => x"02020001",
    23439 => x"00016fbc", 23440 => x"0000c2a0", 23441 => x"00000000",
    23442 => x"00018f34", 23443 => x"02040010", 23444 => x"00016fc0",
    23445 => x"0000c2a0", 23446 => x"00000000", 23447 => x"00018ed0",
    23448 => x"02020004", 23449 => x"00016fc4", 23450 => x"0000c2a0",
    23451 => x"00000000", 23452 => x"0001927c", 23453 => x"02410004",
    23454 => x"00016fc8", 23455 => x"0000c2a0", 23456 => x"00000000",
    23457 => x"00019280", 23458 => x"02410004", 23459 => x"00000000",
    23460 => x"00000000", 23461 => x"00000000", 23462 => x"00000000",
    23463 => x"00000000", 23464 => x"2b060104", 23465 => x"01606501",
    23466 => x"08010000", 23467 => x"00016fcc", 23468 => x"0000bfb8",
    23469 => x"00000000", 23470 => x"00000000", 23471 => x"01040001",
    23472 => x"00016fd0", 23473 => x"0000bfb8", 23474 => x"00000000",
    23475 => x"00000000", 23476 => x"01020001", 23477 => x"00016fd4",
    23478 => x"0000bfb8", 23479 => x"00000000", 23480 => x"00000000",
    23481 => x"01020001", 23482 => x"00016fd8", 23483 => x"0000bfb8",
    23484 => x"00000000", 23485 => x"00000000", 23486 => x"01020001",
    23487 => x"00000000", 23488 => x"00000000", 23489 => x"00000000",
    23490 => x"00000000", 23491 => x"00000000", 23492 => x"01000000",
    23493 => x"02000000", 23494 => x"03000000", 23495 => x"04000000",
    23496 => x"00015608", 23497 => x"01000000", 23498 => x"02000000",
    23499 => x"03000000", 23500 => x"02000000", 23501 => x"03000000",
    23502 => x"01000000", 23503 => x"02000000", 23504 => x"03000000",
    23505 => x"04000000", 23506 => x"05000000", 23507 => x"06000000",
    23508 => x"07000000", 23509 => x"08000000", 23510 => x"09000000",
    23511 => x"05000000", 23512 => x"08000000", 23513 => x"09000000",
    23514 => x"0a000000", 23515 => x"0c000000", 23516 => x"0d000000",
    23517 => x"0e000000", 23518 => x"0f000000", 23519 => x"10000000",
    23520 => x"11000000", 23521 => x"12000000", 23522 => x"13000000",
    23523 => x"14000000", 23524 => x"16000000", 23525 => x"17000000",
    23526 => x"18000000", 23527 => x"1a000000", 23528 => x"01000000",
    23529 => x"02000000", 23530 => x"03000000", 23531 => x"04000000",
    23532 => x"05000000", 23533 => x"06000000", 23534 => x"01000000",
    23535 => x"02000000", 23536 => x"03000000", 23537 => x"04000000",
    23538 => x"05000000", 23539 => x"02000000", 23540 => x"03000000",
    23541 => x"04000000", 23542 => x"05000000", 23543 => x"000171c8",
    23544 => x"000172b4", 23545 => x"00000000", 23546 => x"00000000",
    23547 => x"00000004", 23548 => x"00000008", 23549 => x"00000100",
    23550 => x"00000200", 23551 => x"046362a0", 23552 => x"000192bc",
    23553 => x"00000000", 23554 => x"00000000", 23555 => x"0000ce42",
    23556 => x"ab28633a", 23557 => x"00000000", 23558 => x"00018f28",
    23559 => x"00000000", 23560 => x"00000000", 23561 => x"0000ce42",
    23562 => x"650c2d4f", 23563 => x"00000000", 23564 => x"000192c4",
    23565 => x"00000000", 23566 => x"00000000", 23567 => x"0000ce42",
    23568 => x"65158dc0", 23569 => x"00000000", 23570 => x"00018f48",
    23571 => x"00000000", 23572 => x"00000000", 23573 => x"0000ce42",
    23574 => x"de0d8ced", 23575 => x"00000000", 23576 => x"000192c0",
    23577 => x"00000000", 23578 => x"00000000", 23579 => x"0000ce42",
    23580 => x"ff07fc47", 23581 => x"00000000", 23582 => x"00019288",
    23583 => x"00000000", 23584 => x"00000000", 23585 => x"0000ce42",
    23586 => x"e2d13d04", 23587 => x"00000000", 23588 => x"00019258",
    23589 => x"00000000", 23590 => x"00000000", 23591 => x"0000ce42",
    23592 => x"779c5443", 23593 => x"00000000", 23594 => x"000192b8",
    23595 => x"00000000", 23596 => x"00000000", 23597 => x"00000651",
    23598 => x"68202b22", 23599 => x"00000000", 23600 => x"000192b0",
    23601 => x"00000000", 23602 => x"00000000", 23603 => x"00001103",
    23604 => x"c0413599", 23605 => x"00000000", 23606 => x"0001929c",
    23607 => x"00000000", 23608 => x"00000000", 23609 => x"00001103",
    23610 => x"f0f43591", 23611 => x"00000000", 23612 => x"00015740",
    23613 => x"00000000", 23614 => x"00000001", 23615 => x"00030000",
    23616 => x"00000004", 23617 => x"00000000", 23618 => x"00000000",
    23619 => x"00000000", 23620 => x"00000000", 23621 => x"00000000",
    23622 => x"00000000", 23623 => x"00000000", 23624 => x"00000000",
    23625 => x"00000000", 23626 => x"00000000", 23627 => x"00000000",
    23628 => x"00000000", 23629 => x"00000000", 23630 => x"00000000",
    23631 => x"00000000", 23632 => x"00000000", 23633 => x"00000000",
    23634 => x"00000000", 23635 => x"00000000", 23636 => x"00000000",
    23637 => x"00000000", 23638 => x"00000000", 23639 => x"00000000",
    23640 => x"00000000", 23641 => x"00000000", 23642 => x"00000000",
    23643 => x"00000000", 23644 => x"00000000", 23645 => x"00000000",
    23646 => x"00000000", 23647 => x"00000000", 23648 => x"00000000",
    23649 => x"00000000", 23650 => x"00000000", 23651 => x"00000000",
    23652 => x"00000000", 23653 => x"00000000", 23654 => x"00000000",
    23655 => x"00000000", 23656 => x"00000000", 23657 => x"00000000",
    23658 => x"ff000000", 23659 => x"0000fe50", 23660 => x"0000fe84",
    23661 => x"0000feb4", 23662 => x"00014a80", 23663 => x"80000000",
    23664 => x"00000000", 23665 => x"00000000", 23666 => x"44332211",
    23667 => x"00000000", 23668 => x"04000000", 23669 => x"138046e2",
    23670 => x"01000000", 23671 => x"9000cfea", 23672 => x"01000000",
    23673 => x"108157f3", 23674 => x"01000000", 23675 => x"0be0ffff",
    23676 => x"01000000", 23677 => x"88e0ffff", 23678 => x"01000000",
    23679 => x"08e1ffff", 23680 => x"01000000", 23681 => x"1b0020e0",
    23682 => x"01000000", 23683 => x"9800c0eb", 23684 => x"01000000",
    23685 => x"6b2130e0", 23686 => x"01000000", 23687 => x"69610de0",
    23688 => x"01000000", 23689 => x"10a38900", 23690 => x"04000000",
    23691 => x"33e31ef1", 23692 => x"01000000", 23693 => x"31c35ff9",
    23694 => x"01000000", 23695 => x"2b0300e1", 23696 => x"01000000",
    23697 => x"43c300e1", 23698 => x"01000000", 23699 => x"79411400",
    23700 => x"04000000", 23701 => x"cb250060", 23702 => x"00000000",
    23703 => x"81c88001", 23704 => x"04000000", 23705 => x"c02fc100",
    23706 => x"04000000", 23707 => x"d3250260", 23708 => x"00000000",
    23709 => x"50ea8101", 23710 => x"04000000", 23711 => x"5b090080",
    23712 => x"01000000", 23713 => x"59092080", 23714 => x"01000000",
    23715 => x"c86a8101", 23716 => x"04000000", 23717 => x"63097afd",
    23718 => x"01000000", 23719 => x"e88a8101", 23720 => x"04000000",
    23721 => x"fc8a8101", 23722 => x"04000000", 23723 => x"00000000",
    23724 => x"08000000", 23725 => x"ffffffff", 23726 => x"00016054",
    23727 => x"5b1157a7", 23728 => x"00000003", 23729 => x"00000000",
    23730 => x"00000000", 23731 => x"00000000", 23732 => x"00000000",
    23733 => x"00000000", 23734 => x"00000000", 23735 => x"00000000",
    23736 => x"00000000", 23737 => x"00000000", 23738 => x"00000000",
    23739 => x"00000000", 23740 => x"77727063", 23741 => x"2d76332e",
    23742 => x"302d3238", 23743 => x"322d6763", 23744 => x"35373161",
    23745 => x"31662d64", 23746 => x"69727479", 23747 => x"00000000",
    23748 => x"44656320", 23749 => x"20362032", 23750 => x"30313600",
    23751 => x"00000000", 23752 => x"31303a33", 23753 => x"343a3133",
    23754 => x"00000000", 23755 => x"00000000", 23756 => x"686f6e67",
    23757 => x"6d696e67", 23758 => x"00000000", 23759 => x"00000000",
    23760 => x"00000000", 23761 => x"00000000", 23762 => x"00000000",
    23763 => x"00000000", 23764 => x"00014f90", 23765 => x"00008880",
    23766 => x"0001375c", 23767 => x"00008940", 23768 => x"00014fa8",
    23769 => x"000089a0", 23770 => x"00014fdc", 23771 => x"00008a3c",
    23772 => x"00015030", 23773 => x"00008b54", 23774 => x"00015080",
    23775 => x"00008c64", 23776 => x"000150a0", 23777 => x"00008d44",
    23778 => x"000150c4", 23779 => x"00008da4", 23780 => x"000151f4",
    23781 => x"00008ea8", 23782 => x"00015230", 23783 => x"00009240",
    23784 => x"0001528c", 23785 => x"000094a8", 23786 => x"000152c4",
    23787 => x"00009580", 23788 => x"000152cc", 23789 => x"000096e0",
    23790 => x"000152d0", 23791 => x"000096f8", 23792 => x"00015300",
    23793 => x"00009714", 23794 => x"00015314", 23795 => x"000097c0",
    23796 => x"00015384", 23797 => x"000098e0", 23798 => x"000153a0",
    23799 => x"000099d0", 23800 => x"00015428", 23801 => x"00009a90",
    23802 => x"00015430", 23803 => x"00009a18", 23804 => x"000151f8",
    23805 => x"00009b5c", 23806 => x"00015824", 23807 => x"0000eb94",
    23808 => x"00015938", 23809 => x"00010100", 23810 => x"0001593c",
    23811 => x"00010004", 23812 => x"00015940", 23813 => x"0000ff08",
    23814 => x"00010734", 23815 => x"00000000", 23816 => x"000171b8",
    23817 => x"00013774", 23818 => x"00000000", 23819 => x"00000214",
    23820 => x"00000000", 23821 => x"00000000", 23822 => x"00000000",
    23823 => x"00000000", 23824 => x"00013748", 23825 => x"00000000",
    23826 => x"00000000", 23827 => x"00012450", 23828 => x"00000000",
    23829 => x"00000000", 23830 => x"00000000", 23831 => x"00013750",
    23832 => x"00000000", 23833 => x"000087d4", 23834 => x"000004f8",
    23835 => x"00000000", 23836 => x"00000000", 23837 => x"00000000",
    23838 => x"0001375c", 23839 => x"00000000", 23840 => x"00000000",
    23841 => x"000010e8", 23842 => x"00000000", 23843 => x"00000000",
    23844 => x"00000000", 23845 => x"00013760", 23846 => x"00000000",
    23847 => x"000004d4", 23848 => x"00000468", 23849 => x"00000000",
    23850 => x"00000000", 23851 => x"00000000", 23852 => x"00013768",
    23853 => x"00000000", 23854 => x"00000000", 23855 => x"00000378",
    23856 => x"00000000", 23857 => x"00000000", 23858 => x"00000000",
    23859 => x"00014e78", 23860 => x"00000000", 23861 => x"00000000",
    23862 => x"00007678", 23863 => x"00000000", 23864 => x"00000000",
    23865 => x"00000000", 23866 => x"00015588", 23867 => x"000192a0",
    23868 => x"00000000", 23869 => x"0000a298", 23870 => x"00000000",
    23871 => x"00000000", 23872 => x"00000000", 23873 => x"00015590",
    23874 => x"000192a0", 23875 => x"0000aa08", 23876 => x"0000aab8",
    23877 => x"00000000", 23878 => x"00000000", 23879 => x"00000000",
    23880 => x"00015598", 23881 => x"000192a0", 23882 => x"0000afc4",
    23883 => x"0000ae38", 23884 => x"00000000", 23885 => x"00000000",
    23886 => x"00000000", 23887 => x"00015600", 23888 => x"000192a0",
    23889 => x"0000c6e4", 23890 => x"0000b70c", 23891 => x"00000000",
    23892 => x"00000000", 23893 => x"00000000", 23894 => x"0001582c",
    23895 => x"00000000", 23896 => x"0000e86c", 23897 => x"0000e8b8",
    23898 => x"00000000", 23899 => x"00000000", 23900 => x"00000000",
    23901 => x"00000000", 23902 => x"00000000", 23903 => x"00000000",
    23904 => x"00000000", 23905 => x"00000000", 23906 => x"00000000",
    23907 => x"00000000", 23908 => x"00000000", 23909 => x"00000000",
    23910 => x"00000000", 23911 => x"00000000", 23912 => x"00000000",
    23913 => x"00000000", 23914 => x"00000000", 23915 => x"00000000",
    23916 => x"00000000", 23917 => x"00000000", 23918 => x"00000000",
    23919 => x"00000000", 23920 => x"00000000", 23921 => x"00000000",
    23922 => x"00000000", 23923 => x"00000000", 23924 => x"00000000",
    23925 => x"00000000", 23926 => x"00000000", 23927 => x"00000000",
    23928 => x"00000000", 23929 => x"00000000", 23930 => x"00000000",
    23931 => x"00000000", 23932 => x"00000000", 23933 => x"00000000",
    23934 => x"00000000", 23935 => x"00000000", 23936 => x"00000000",
    23937 => x"00000000", 23938 => x"00000000", 23939 => x"00000000",
    23940 => x"00000000", 23941 => x"00000000", 23942 => x"00000000",
    23943 => x"00000000", 23944 => x"00000000", 23945 => x"00000000",
    23946 => x"00000000", 23947 => x"00000000", 23948 => x"00000000",
    23949 => x"00000000", 23950 => x"00000000", 23951 => x"00000000",
    23952 => x"00000000", 23953 => x"00000000", 23954 => x"00000000",
    23955 => x"00000000", 23956 => x"00000000", 23957 => x"00000000",
    23958 => x"00000000", 23959 => x"00000000", 23960 => x"00000000",
    23961 => x"00000000", 23962 => x"00000000", 23963 => x"00000000",
    23964 => x"00000000", 23965 => x"00000000", 23966 => x"00000000",
    23967 => x"00000000", 23968 => x"00000000", 23969 => x"00000000",
    23970 => x"00000000", 23971 => x"00000000", 23972 => x"00000000",
    23973 => x"00000000", 23974 => x"00000000", 23975 => x"00000000",
    23976 => x"00000000", 23977 => x"00000000", 23978 => x"00000000",
    23979 => x"00000000", 23980 => x"00000000", 23981 => x"00000000",
    23982 => x"00000000", 23983 => x"00000000", 23984 => x"00000000",
    23985 => x"00000000", 23986 => x"00000000", 23987 => x"00000000",
    23988 => x"00000000", 23989 => x"00000000", 23990 => x"00000000",
    23991 => x"00000000", 23992 => x"00000000", 23993 => x"00000000",
    23994 => x"00000000", 23995 => x"00000000", 23996 => x"00000000",
    23997 => x"00000000", 23998 => x"00000000", 23999 => x"00000000",
    24000 => x"00000000", 24001 => x"00000000", 24002 => x"00000000",
    24003 => x"00000000", 24004 => x"00000000", 24005 => x"00000000",
    24006 => x"00000000", 24007 => x"00000000", 24008 => x"00000000",
    24009 => x"00000000", 24010 => x"00000000", 24011 => x"00000000",
    24012 => x"00000000", 24013 => x"00000000", 24014 => x"00000000",
    24015 => x"00000000", 24016 => x"00000000", 24017 => x"00000000",
    24018 => x"00000000", 24019 => x"00000000", 24020 => x"00000000",
    24021 => x"00000000", 24022 => x"00000000", 24023 => x"00000000",
    24024 => x"00000000", 24025 => x"00000000", 24026 => x"00000000",
    24027 => x"00000000", 24028 => x"00000000", 24029 => x"00000000",
    24030 => x"00000000", 24031 => x"00000000", 24032 => x"00000000",
    24033 => x"00000000", 24034 => x"00000000", 24035 => x"00000000",
    24036 => x"00000000", 24037 => x"00000000", 24038 => x"00000000",
    24039 => x"00000000", 24040 => x"00000000", 24041 => x"00000000",
    24042 => x"00000000", 24043 => x"00000000", 24044 => x"00000000",
    24045 => x"00000000", 24046 => x"00000000", 24047 => x"00000000",
    24048 => x"00000000", 24049 => x"00000000", 24050 => x"00000000",
    24051 => x"00000000", 24052 => x"00000000", 24053 => x"00000000",
    24054 => x"00000000", 24055 => x"00000000", 24056 => x"00000000",
    24057 => x"00000000", 24058 => x"00000000", 24059 => x"00000000",
    24060 => x"00000000", 24061 => x"00000000", 24062 => x"00000000",
    24063 => x"00000000", 24064 => x"00000000", 24065 => x"00000000",
    24066 => x"00000000", 24067 => x"00000000", 24068 => x"00000000",
    24069 => x"00000000", 24070 => x"00000000", 24071 => x"00000000",
    24072 => x"00000000", 24073 => x"00000000", 24074 => x"00000000",
    24075 => x"00000000", 24076 => x"00000000", 24077 => x"00000000",
    24078 => x"00000000", 24079 => x"00000000", 24080 => x"00000000",
    24081 => x"00000000", 24082 => x"00000000", 24083 => x"00000000",
    24084 => x"00000000", 24085 => x"00000000", 24086 => x"00000000",
    24087 => x"00000000", 24088 => x"00000000", 24089 => x"00000000",
    24090 => x"00000000", 24091 => x"00000000", 24092 => x"00000000",
    24093 => x"00000000", 24094 => x"00000000", 24095 => x"00000000",
    24096 => x"00000000", 24097 => x"00000000", 24098 => x"00000000",
    24099 => x"00000000", 24100 => x"00000000", 24101 => x"00000000",
    24102 => x"00000000", 24103 => x"00000000", 24104 => x"00000000",
    24105 => x"00000000", 24106 => x"00000000", 24107 => x"00000000",
    24108 => x"00000000", 24109 => x"00000000", 24110 => x"00000000",
    24111 => x"00000000", 24112 => x"00000000", 24113 => x"00000000",
    24114 => x"00000000", 24115 => x"00000000", 24116 => x"00000000",
    24117 => x"00000000", 24118 => x"00000000", 24119 => x"00000000",
    24120 => x"00000000", 24121 => x"00000000", 24122 => x"00000000",
    24123 => x"00000000", 24124 => x"00000000", 24125 => x"00000000",
    24126 => x"00000000", 24127 => x"00000000", 24128 => x"00000000",
    24129 => x"00000000", 24130 => x"00000000", 24131 => x"00000000",
    24132 => x"00000000", 24133 => x"00000000", 24134 => x"00000000",
    24135 => x"00000000", 24136 => x"00000000", 24137 => x"00000000",
    24138 => x"00000000", 24139 => x"00000000", 24140 => x"00000000",
    24141 => x"00000000", 24142 => x"00000000", 24143 => x"00000000",
    24144 => x"00000000", 24145 => x"00000000", 24146 => x"00000000",
    24147 => x"00000000", 24148 => x"00000000", 24149 => x"00000000",
    24150 => x"00000000", 24151 => x"00000000", 24152 => x"00000000",
    24153 => x"00000000", 24154 => x"00000000", 24155 => x"00000000",
    24156 => x"00000000", 24157 => x"00000000", 24158 => x"00000000",
    24159 => x"00000000", 24160 => x"00000000", 24161 => x"00000000",
    24162 => x"00000000", 24163 => x"00000000", 24164 => x"00000000",
    24165 => x"00000000", 24166 => x"00000000", 24167 => x"00000000",
    24168 => x"00000000", 24169 => x"00000000", 24170 => x"00000000",
    24171 => x"00000000", 24172 => x"00000000", 24173 => x"00000000",
    24174 => x"00000000", 24175 => x"00000000", 24176 => x"00000000",
    24177 => x"00000000", 24178 => x"00000000", 24179 => x"00000000",
    24180 => x"00000000", 24181 => x"00000000", 24182 => x"00000000",
    24183 => x"00000000", 24184 => x"00000000", 24185 => x"00000000",
    24186 => x"00000000", 24187 => x"00000000", 24188 => x"00000000",
    24189 => x"00000000", 24190 => x"00000000", 24191 => x"00000000",
    24192 => x"00000000", 24193 => x"00000000", 24194 => x"00000000",
    24195 => x"00000000", 24196 => x"00000000", 24197 => x"00000000",
    24198 => x"00000000", 24199 => x"00000000", 24200 => x"00000000",
    24201 => x"00000000", 24202 => x"00000000", 24203 => x"00000000",
    24204 => x"00000000", 24205 => x"00000000", 24206 => x"00000000",
    24207 => x"00000000", 24208 => x"00000000", 24209 => x"00000000",
    24210 => x"00000000", 24211 => x"00000000", 24212 => x"00000000",
    24213 => x"00000000", 24214 => x"00000000", 24215 => x"00000000",
    24216 => x"00000000", 24217 => x"00000000", 24218 => x"00000000",
    24219 => x"00000000", 24220 => x"00000000", 24221 => x"00000000",
    24222 => x"00000000", 24223 => x"00000000", 24224 => x"00000000",
    24225 => x"00000000", 24226 => x"00000000", 24227 => x"00000000",
    24228 => x"00000000", 24229 => x"00000000", 24230 => x"00000000",
    24231 => x"00000000", 24232 => x"00000000", 24233 => x"00000000",
    24234 => x"00000000", 24235 => x"00000000", 24236 => x"00000000",
    24237 => x"00000000", 24238 => x"00000000", 24239 => x"00000000",
    24240 => x"00000000", 24241 => x"00000000", 24242 => x"00000000",
    24243 => x"00000000", 24244 => x"00000000", 24245 => x"00000000",
    24246 => x"00000000", 24247 => x"00000000", 24248 => x"00000000",
    24249 => x"00000000", 24250 => x"00000000", 24251 => x"00000000",
    24252 => x"00000000", 24253 => x"00000000", 24254 => x"00000000",
    24255 => x"00000000", 24256 => x"00000000", 24257 => x"00000000",
    24258 => x"00000000", 24259 => x"00000000", 24260 => x"00000000",
    24261 => x"00000000", 24262 => x"00000000", 24263 => x"00000000",
    24264 => x"00000000", 24265 => x"00000000", 24266 => x"00000000",
    24267 => x"00000000", 24268 => x"00000000", 24269 => x"00000000",
    24270 => x"00000000", 24271 => x"00000000", 24272 => x"00000000",
    24273 => x"00000000", 24274 => x"00000000", 24275 => x"00000000",
    24276 => x"00000000", 24277 => x"00000000", 24278 => x"00000000",
    24279 => x"00000000", 24280 => x"00000000", 24281 => x"00000000",
    24282 => x"00000000", 24283 => x"00000000", 24284 => x"00000000",
    24285 => x"00000000", 24286 => x"00000000", 24287 => x"00000000",
    24288 => x"00000000", 24289 => x"00000000", 24290 => x"00000000",
    24291 => x"00000000", 24292 => x"00000000", 24293 => x"00000000",
    24294 => x"00000000", 24295 => x"00000000", 24296 => x"00000000",
    24297 => x"00000000", 24298 => x"00000000", 24299 => x"00000000",
    24300 => x"00000000", 24301 => x"00000000", 24302 => x"00000000",
    24303 => x"00000000", 24304 => x"00000000", 24305 => x"00000000",
    24306 => x"00000000", 24307 => x"00000000", 24308 => x"00000000",
    24309 => x"00000000", 24310 => x"00000000", 24311 => x"00000000",
    24312 => x"00000000", 24313 => x"00000000", 24314 => x"00000000",
    24315 => x"00000000", 24316 => x"00000000", 24317 => x"00000000",
    24318 => x"00000000", 24319 => x"00000000", 24320 => x"00000000",
    24321 => x"00000000", 24322 => x"00000000", 24323 => x"00000000",
    24324 => x"00000000", 24325 => x"00000000", 24326 => x"00000000",
    24327 => x"00000000", 24328 => x"00000000", 24329 => x"00000000",
    24330 => x"00000000", 24331 => x"00000000", 24332 => x"00000000",
    24333 => x"00000000", 24334 => x"00000000", 24335 => x"00000000",
    24336 => x"00000000", 24337 => x"00000000", 24338 => x"00000000",
    24339 => x"00000000", 24340 => x"00000000", 24341 => x"00000000",
    24342 => x"00000000", 24343 => x"00000000", 24344 => x"00000000",
    24345 => x"00000000", 24346 => x"00000000", 24347 => x"00000000",
    24348 => x"00000000", 24349 => x"00000000", 24350 => x"00000000",
    24351 => x"00000000", 24352 => x"00000000", 24353 => x"00000000",
    24354 => x"00000000", 24355 => x"00000000", 24356 => x"00000000",
    24357 => x"00000000", 24358 => x"00000000", 24359 => x"00000000",
    24360 => x"00000000", 24361 => x"00000000", 24362 => x"00000000",
    24363 => x"00000000", 24364 => x"00000000", 24365 => x"00000000",
    24366 => x"00000000", 24367 => x"00000000", 24368 => x"00000000",
    24369 => x"00000000", 24370 => x"00000000", 24371 => x"00000000",
    24372 => x"00000000", 24373 => x"00000000", 24374 => x"00000000",
    24375 => x"00000000", 24376 => x"00000000", 24377 => x"00000000",
    24378 => x"00000000", 24379 => x"00000000", 24380 => x"00000000",
    24381 => x"00000000", 24382 => x"00000000", 24383 => x"00000000",
    24384 => x"00000000", 24385 => x"00000000", 24386 => x"00000000",
    24387 => x"00000000", 24388 => x"00000000", 24389 => x"00000000",
    24390 => x"00000000", 24391 => x"00000000", 24392 => x"00000000",
    24393 => x"00000000", 24394 => x"00000000", 24395 => x"00000000",
    24396 => x"00000000", 24397 => x"00000000", 24398 => x"00000000",
    24399 => x"00000000", 24400 => x"00000000", 24401 => x"00000000",
    24402 => x"00000000", 24403 => x"00000000", 24404 => x"00000000",
    24405 => x"00000000", 24406 => x"00000000", 24407 => x"00000000",
    24408 => x"00000000", 24409 => x"00000000", 24410 => x"00000000",
    24411 => x"00000000", 24412 => x"00000000", 24413 => x"00000000",
    24414 => x"00000000", 24415 => x"00000000", 24416 => x"00000000",
    24417 => x"00000000", 24418 => x"00000000", 24419 => x"00000000",
    24420 => x"00000000", 24421 => x"00000000", 24422 => x"00000000",
    24423 => x"00000000", 24424 => x"00000000", 24425 => x"00000000",
    24426 => x"00000000", 24427 => x"00000000", 24428 => x"00000000",
    24429 => x"00000000", 24430 => x"00000000", 24431 => x"00000000",
    24432 => x"00000000", 24433 => x"00000000", 24434 => x"00000000",
    24435 => x"00000000", 24436 => x"00000000", 24437 => x"00000000",
    24438 => x"00000000", 24439 => x"00000000", 24440 => x"00000000",
    24441 => x"00000000", 24442 => x"00000000", 24443 => x"00000000",
    24444 => x"00000000", 24445 => x"00000000", 24446 => x"00000000",
    24447 => x"00000000", 24448 => x"00000000", 24449 => x"00000000",
    24450 => x"00000000", 24451 => x"00000000", 24452 => x"00000000",
    24453 => x"00000000", 24454 => x"00000000", 24455 => x"00000000",
    24456 => x"00000000", 24457 => x"00000000", 24458 => x"00000000",
    24459 => x"00000000", 24460 => x"00000000", 24461 => x"00000000",
    24462 => x"00000000", 24463 => x"00000000", 24464 => x"00000000",
    24465 => x"00000000", 24466 => x"00000000", 24467 => x"00000000",
    24468 => x"00000000", 24469 => x"00000000", 24470 => x"00000000",
    24471 => x"00000000", 24472 => x"00000000", 24473 => x"00000000",
    24474 => x"00000000", 24475 => x"00000000", 24476 => x"00000000",
    24477 => x"00000000", 24478 => x"00000000", 24479 => x"00000000",
    24480 => x"00000000", 24481 => x"00000000", 24482 => x"00000000",
    24483 => x"00000000", 24484 => x"00000000", 24485 => x"00000000",
    24486 => x"00000000", 24487 => x"00000000", 24488 => x"00000000",
    24489 => x"00000000", 24490 => x"00000000", 24491 => x"00000000",
    24492 => x"00000000", 24493 => x"00000000", 24494 => x"00000000",
    24495 => x"00000000", 24496 => x"00000000", 24497 => x"00000000",
    24498 => x"00000000", 24499 => x"00000000", 24500 => x"00000000",
    24501 => x"00000000", 24502 => x"00000000", 24503 => x"00000000",
    24504 => x"00000000", 24505 => x"00000000", 24506 => x"00000000",
    24507 => x"00000000", 24508 => x"00000000", 24509 => x"00000000",
    24510 => x"00000000", 24511 => x"00000000", 24512 => x"00000000",
    24513 => x"00000000", 24514 => x"00000000", 24515 => x"00000000",
    24516 => x"00000000", 24517 => x"00000000", 24518 => x"00000000",
    24519 => x"00000000", 24520 => x"00000000", 24521 => x"00000000",
    24522 => x"00000000", 24523 => x"00000000", 24524 => x"00000000",
    24525 => x"00000000", 24526 => x"00000000", 24527 => x"00000000",
    24528 => x"00000000", 24529 => x"00000000", 24530 => x"00000000",
    24531 => x"00000000", 24532 => x"00000000", 24533 => x"00000000",
    24534 => x"00000000", 24535 => x"00000000", 24536 => x"00000000",
    24537 => x"00000000", 24538 => x"00000000", 24539 => x"00000000",
    24540 => x"00000000", 24541 => x"00000000", 24542 => x"00000000",
    24543 => x"00000000", 24544 => x"00000000", 24545 => x"00000000",
    24546 => x"00000000", 24547 => x"00000000", 24548 => x"00000000",
    24549 => x"00000000", 24550 => x"00000000", 24551 => x"00000000",
    24552 => x"00000000", 24553 => x"00000000", 24554 => x"00000000",
    24555 => x"00000000", 24556 => x"00000000", 24557 => x"00000000",
    24558 => x"00000000", 24559 => x"00000000", 24560 => x"00000000",
    24561 => x"00000000", 24562 => x"00000000", 24563 => x"00000000",
    24564 => x"00000000", 24565 => x"00000000", 24566 => x"00000000",
    24567 => x"00000000", 24568 => x"00000000", 24569 => x"00000000",
    24570 => x"00000000", 24571 => x"00000000", 24572 => x"00000000",
    24573 => x"00000000", 24574 => x"00000000", 24575 => x"00000000",
    24576 => x"00000000", 24577 => x"00000000", 24578 => x"00000000",
    24579 => x"00000000", 24580 => x"00000000", 24581 => x"00000000",
    24582 => x"00000000", 24583 => x"00000000", 24584 => x"00000000",
    24585 => x"00000000", 24586 => x"00000000", 24587 => x"00000000",
    24588 => x"00000000", 24589 => x"00000000", 24590 => x"00000000",
    24591 => x"00000000", 24592 => x"00000000", 24593 => x"00000000",
    24594 => x"00000000", 24595 => x"00000000", 24596 => x"00000000",
    24597 => x"00000000", 24598 => x"00000000", 24599 => x"00000000",
    24600 => x"00000000", 24601 => x"00000000", 24602 => x"00000000",
    24603 => x"00000000", 24604 => x"00000000", 24605 => x"00000000",
    24606 => x"00000000", 24607 => x"00000000", 24608 => x"00000000",
    24609 => x"00000000", 24610 => x"00000000", 24611 => x"00000000",
    24612 => x"00000000", 24613 => x"00000000", 24614 => x"00000000",
    24615 => x"00000000", 24616 => x"00000000", 24617 => x"00000000",
    24618 => x"00000000", 24619 => x"00000000", 24620 => x"00000000",
    24621 => x"00000000", 24622 => x"00000000", 24623 => x"00000000",
    24624 => x"00000000", 24625 => x"00000000", 24626 => x"00000000",
    24627 => x"00000000", 24628 => x"00000000", 24629 => x"00000000",
    24630 => x"00000000", 24631 => x"00000000", 24632 => x"00000000",
    24633 => x"00000000", 24634 => x"00000000", 24635 => x"00000000",
    24636 => x"00000000", 24637 => x"00000000", 24638 => x"00000000",
    24639 => x"00000000", 24640 => x"00000000", 24641 => x"00000000",
    24642 => x"00000000", 24643 => x"00000000", 24644 => x"00000000",
    24645 => x"00000000", 24646 => x"00000000", 24647 => x"00000000",
    24648 => x"00000000", 24649 => x"00000000", 24650 => x"00000000",
    24651 => x"00000000", 24652 => x"00000000", 24653 => x"00000000",
    24654 => x"00000000", 24655 => x"00000000", 24656 => x"00000000",
    24657 => x"00000000", 24658 => x"00000000", 24659 => x"00000000",
    24660 => x"00000000", 24661 => x"00000000", 24662 => x"00000000",
    24663 => x"00000000", 24664 => x"00000000", 24665 => x"00000000",
    24666 => x"00000000", 24667 => x"00000000", 24668 => x"00000000",
    24669 => x"00000000", 24670 => x"00000000", 24671 => x"00000000",
    24672 => x"00000000", 24673 => x"00000000", 24674 => x"00000000",
    24675 => x"00000000", 24676 => x"00000000", 24677 => x"00000000",
    24678 => x"00000000", 24679 => x"00000000", 24680 => x"00000000",
    24681 => x"00000000", 24682 => x"00000000", 24683 => x"00000000",
    24684 => x"00000000", 24685 => x"00000000", 24686 => x"00000000",
    24687 => x"00000000", 24688 => x"00000000", 24689 => x"00000000",
    24690 => x"00000000", 24691 => x"00000000", 24692 => x"00000000",
    24693 => x"00000000", 24694 => x"00000000", 24695 => x"00000000",
    24696 => x"00000000", 24697 => x"00000000", 24698 => x"00000000",
    24699 => x"00000000", 24700 => x"00000000", 24701 => x"00000000",
    24702 => x"00000000", 24703 => x"00000000", 24704 => x"00000000",
    24705 => x"00000000", 24706 => x"00000000", 24707 => x"00000000",
    24708 => x"00000000", 24709 => x"00000000", 24710 => x"00000000",
    24711 => x"00000000", 24712 => x"00000000", 24713 => x"00000000",
    24714 => x"00000000", 24715 => x"00000000", 24716 => x"00000000",
    24717 => x"00000000", 24718 => x"00000000", 24719 => x"00000000",
    24720 => x"00000000", 24721 => x"00000000", 24722 => x"00000000",
    24723 => x"00000000", 24724 => x"00000000", 24725 => x"00000000",
    24726 => x"00000000", 24727 => x"00000000", 24728 => x"00000000",
    24729 => x"00000000", 24730 => x"00000000", 24731 => x"00000000",
    24732 => x"00000000", 24733 => x"00000000", 24734 => x"00000000",
    24735 => x"00000000", 24736 => x"00000000", 24737 => x"00000000",
    24738 => x"00000000", 24739 => x"00000000", 24740 => x"00000000",
    24741 => x"00000000", 24742 => x"00000000", 24743 => x"00000000",
    24744 => x"00000000", 24745 => x"00000000", 24746 => x"00000000",
    24747 => x"00000000", 24748 => x"00000000", 24749 => x"00000000",
    24750 => x"00000000", 24751 => x"00000000", 24752 => x"00000000",
    24753 => x"00000000", 24754 => x"00000000", 24755 => x"00000000",
    24756 => x"00000000", 24757 => x"00000000", 24758 => x"00000000",
    24759 => x"00000000", 24760 => x"00000000", 24761 => x"00000000",
    24762 => x"00000000", 24763 => x"00000000", 24764 => x"00000000",
    24765 => x"00000000", 24766 => x"00000000", 24767 => x"00000000",
    24768 => x"00000000", 24769 => x"00000000", 24770 => x"00000000",
    24771 => x"00000000", 24772 => x"00000000", 24773 => x"00000000",
    24774 => x"00000000", 24775 => x"00000000", 24776 => x"00000000",
    24777 => x"00000000", 24778 => x"00000000", 24779 => x"00000000",
    24780 => x"00000000", 24781 => x"00000000", 24782 => x"00000000",
    24783 => x"00000000", 24784 => x"00000000", 24785 => x"00000000",
    24786 => x"00000000", 24787 => x"00000000", 24788 => x"00000000",
    24789 => x"00000000", 24790 => x"00000000", 24791 => x"00000000",
    24792 => x"00000000", 24793 => x"00000000", 24794 => x"00000000",
    24795 => x"00000000", 24796 => x"00000000", 24797 => x"00000000",
    24798 => x"00000000", 24799 => x"00000000", 24800 => x"00000000",
    24801 => x"00000000", 24802 => x"00000000", 24803 => x"00000000",
    24804 => x"00000000", 24805 => x"00000000", 24806 => x"00000000",
    24807 => x"00000000", 24808 => x"00000000", 24809 => x"00000000",
    24810 => x"00000000", 24811 => x"00000000", 24812 => x"00000000",
    24813 => x"00000000", 24814 => x"00000000", 24815 => x"00000000",
    24816 => x"00000000", 24817 => x"00000000", 24818 => x"00000000",
    24819 => x"00000000", 24820 => x"00000000", 24821 => x"00000000",
    24822 => x"00000000", 24823 => x"00000000", 24824 => x"00000000",
    24825 => x"00000000", 24826 => x"00000000", 24827 => x"00000000",
    24828 => x"00000000", 24829 => x"00000000", 24830 => x"00000000",
    24831 => x"00000000", 24832 => x"00000000", 24833 => x"00000000",
    24834 => x"00000000", 24835 => x"00000000", 24836 => x"00000000",
    24837 => x"00000000", 24838 => x"00000000", 24839 => x"00000000",
    24840 => x"00000000", 24841 => x"00000000", 24842 => x"00000000",
    24843 => x"00000000", 24844 => x"00000000", 24845 => x"00000000",
    24846 => x"00000000", 24847 => x"00000000", 24848 => x"00000000",
    24849 => x"00000000", 24850 => x"00000000", 24851 => x"00000000",
    24852 => x"00000000", 24853 => x"00000000", 24854 => x"00000000",
    24855 => x"00000000", 24856 => x"00000000", 24857 => x"00000000",
    24858 => x"00000000", 24859 => x"00000000", 24860 => x"00000000",
    24861 => x"00000000", 24862 => x"00000000", 24863 => x"00000000",
    24864 => x"00000000", 24865 => x"00000000", 24866 => x"00000000",
    24867 => x"00000000", 24868 => x"00000000", 24869 => x"00000000",
    24870 => x"00000000", 24871 => x"00000000", 24872 => x"00000000",
    24873 => x"00000000", 24874 => x"00000000", 24875 => x"00000000",
    24876 => x"00000000", 24877 => x"00000000", 24878 => x"00000000",
    24879 => x"00000000", 24880 => x"00000000", 24881 => x"00000000",
    24882 => x"00000000", 24883 => x"00000000", 24884 => x"00000000",
    24885 => x"00000000", 24886 => x"00000000", 24887 => x"00000000",
    24888 => x"00000000", 24889 => x"00000000", 24890 => x"00000000",
    24891 => x"00000000", 24892 => x"00000000", 24893 => x"00000000",
    24894 => x"00000000", 24895 => x"00000000", 24896 => x"00000000",
    24897 => x"00000000", 24898 => x"00000000", 24899 => x"00000000",
    24900 => x"00000000", 24901 => x"00000000", 24902 => x"00000000",
    24903 => x"00000000", 24904 => x"00000000", 24905 => x"00000000",
    24906 => x"00000000", 24907 => x"00000000", 24908 => x"00000000",
    24909 => x"00000000", 24910 => x"00000000", 24911 => x"00000000",
    24912 => x"00000000", 24913 => x"00000000", 24914 => x"00000000",
    24915 => x"00000000", 24916 => x"00000000", 24917 => x"00000000",
    24918 => x"00000000", 24919 => x"00000000", 24920 => x"00000000",
    24921 => x"00000000", 24922 => x"00000000", 24923 => x"00000000",
    24924 => x"00000000", 24925 => x"00000000", 24926 => x"00000000",
    24927 => x"00000000", 24928 => x"00000000", 24929 => x"00000000",
    24930 => x"00000000", 24931 => x"00000000", 24932 => x"00000000",
    24933 => x"00000000", 24934 => x"00000000", 24935 => x"00000000",
    24936 => x"00000000", 24937 => x"00000000", 24938 => x"00000000",
    24939 => x"00000000", 24940 => x"00000000", 24941 => x"00000000",
    24942 => x"00000000", 24943 => x"00000000", 24944 => x"00000000",
    24945 => x"00000000", 24946 => x"00000000", 24947 => x"00000000",
    24948 => x"00000000", 24949 => x"00000000", 24950 => x"00000000",
    24951 => x"00000000", 24952 => x"00000000", 24953 => x"00000000",
    24954 => x"00000000", 24955 => x"00000000", 24956 => x"00000000",
    24957 => x"00000000", 24958 => x"00000000", 24959 => x"00000000",
    24960 => x"00000000", 24961 => x"00000000", 24962 => x"00000000",
    24963 => x"00000000", 24964 => x"00000000", 24965 => x"00000000",
    24966 => x"00000000", 24967 => x"00000000", 24968 => x"00000000",
    24969 => x"00000000", 24970 => x"00000000", 24971 => x"00000000",
    24972 => x"00000000", 24973 => x"00000000", 24974 => x"00000000",
    24975 => x"00000000", 24976 => x"00000000", 24977 => x"00000000",
    24978 => x"00000000", 24979 => x"00000000", 24980 => x"00000000",
    24981 => x"00000000", 24982 => x"00000000", 24983 => x"00000000",
    24984 => x"00000000", 24985 => x"00000000", 24986 => x"00000000",
    24987 => x"00000000", 24988 => x"00000000", 24989 => x"00000000",
    24990 => x"00000000", 24991 => x"00000000", 24992 => x"00000000",
    24993 => x"00000000", 24994 => x"00000000", 24995 => x"00000000",
    24996 => x"00000000", 24997 => x"00000000", 24998 => x"00000000",
    24999 => x"00000000", 25000 => x"00000000", 25001 => x"00000000",
    25002 => x"00000000", 25003 => x"00000000", 25004 => x"00000000",
    25005 => x"00000000", 25006 => x"00000000", 25007 => x"00000000",
    25008 => x"00000000", 25009 => x"00000000", 25010 => x"00000000",
    25011 => x"00000000", 25012 => x"00000000", 25013 => x"00000000",
    25014 => x"00000000", 25015 => x"00000000", 25016 => x"00000000",
    25017 => x"00000000", 25018 => x"00000000", 25019 => x"00000000",
    25020 => x"00000000", 25021 => x"00000000", 25022 => x"00000000",
    25023 => x"00000000", 25024 => x"00000000", 25025 => x"00000000",
    25026 => x"00000000", 25027 => x"00000000", 25028 => x"00000000",
    25029 => x"00000000", 25030 => x"00000000", 25031 => x"00000000",
    25032 => x"00000000", 25033 => x"00000000", 25034 => x"00000000",
    25035 => x"00000000", 25036 => x"00000000", 25037 => x"00000000",
    25038 => x"00000000", 25039 => x"00000000", 25040 => x"00000000",
    25041 => x"00000000", 25042 => x"00000000", 25043 => x"00000000",
    25044 => x"00000000", 25045 => x"00000000", 25046 => x"00000000",
    25047 => x"00000000", 25048 => x"00000000", 25049 => x"00000000",
    25050 => x"00000000", 25051 => x"00000000", 25052 => x"00000000",
    25053 => x"00000000", 25054 => x"00000000", 25055 => x"00000000",
    25056 => x"00000000", 25057 => x"00000000", 25058 => x"00000000",
    25059 => x"00000000", 25060 => x"00000000", 25061 => x"00000000",
    25062 => x"00000000", 25063 => x"00000000", 25064 => x"00000000",
    25065 => x"00000000", 25066 => x"00000000", 25067 => x"00000000",
    25068 => x"00000000", 25069 => x"00000000", 25070 => x"00000000",
    25071 => x"00000000", 25072 => x"00000000", 25073 => x"00000000",
    25074 => x"00000000", 25075 => x"00000000", 25076 => x"00000000",
    25077 => x"00000000", 25078 => x"00000000", 25079 => x"00000000",
    25080 => x"00000000", 25081 => x"00000000", 25082 => x"00000000",
    25083 => x"00000000", 25084 => x"00000000", 25085 => x"00000000",
    25086 => x"00000000", 25087 => x"00000000", 25088 => x"00000000",
    25089 => x"00000000", 25090 => x"00000000", 25091 => x"00000000",
    25092 => x"00000000", 25093 => x"00000000", 25094 => x"00000000",
    25095 => x"00000000", 25096 => x"00000000", 25097 => x"00000000",
    25098 => x"00000000", 25099 => x"00000000", 25100 => x"00000000",
    25101 => x"00000000", 25102 => x"00000000", 25103 => x"00000000",
    25104 => x"00000000", 25105 => x"00000000", 25106 => x"00000000",
    25107 => x"00000000", 25108 => x"00000000", 25109 => x"00000000",
    25110 => x"00000000", 25111 => x"00000000", 25112 => x"00000000",
    25113 => x"00000000", 25114 => x"00000000", 25115 => x"00000000",
    25116 => x"00000000", 25117 => x"00000000", 25118 => x"00000000",
    25119 => x"00000000", 25120 => x"00000000", 25121 => x"00000000",
    25122 => x"00000000", 25123 => x"00000000", 25124 => x"00000000",
    25125 => x"00000000", 25126 => x"00000000", 25127 => x"00000000",
    25128 => x"00000000", 25129 => x"00000000", 25130 => x"00000000",
    25131 => x"00000000", 25132 => x"00000000", 25133 => x"00000000",
    25134 => x"00000000", 25135 => x"00000000", 25136 => x"00000000",
    25137 => x"00000000", 25138 => x"00000000", 25139 => x"00000000",
    25140 => x"00000000", 25141 => x"00000000", 25142 => x"00000000",
    25143 => x"00000000", 25144 => x"00000000", 25145 => x"00000000",
    25146 => x"00000000", 25147 => x"00000000", 25148 => x"00000000",
    25149 => x"00000000", 25150 => x"00000000", 25151 => x"00000000",
    25152 => x"00000000", 25153 => x"00000000", 25154 => x"00000000",
    25155 => x"00000000", 25156 => x"00000000", 25157 => x"00000000",
    25158 => x"00000000", 25159 => x"00000000", 25160 => x"00000000",
    25161 => x"00000000", 25162 => x"00000000", 25163 => x"00000000",
    25164 => x"00000000", 25165 => x"00000000", 25166 => x"00000000",
    25167 => x"00000000", 25168 => x"00000000", 25169 => x"00000000",
    25170 => x"00000000", 25171 => x"00000000", 25172 => x"00000000",
    25173 => x"00000000", 25174 => x"00000000", 25175 => x"00000000",
    25176 => x"00000000", 25177 => x"00000000", 25178 => x"00000000",
    25179 => x"00000000", 25180 => x"00000000", 25181 => x"00000000",
    25182 => x"00000000", 25183 => x"00000000", 25184 => x"00000000",
    25185 => x"00000000", 25186 => x"00000000", 25187 => x"00000000",
    25188 => x"00000000", 25189 => x"00000000", 25190 => x"00000000",
    25191 => x"00000000", 25192 => x"00000000", 25193 => x"00000000",
    25194 => x"00000000", 25195 => x"00000000", 25196 => x"00000000",
    25197 => x"00000000", 25198 => x"00000000", 25199 => x"00000000",
    25200 => x"00000000", 25201 => x"00000000", 25202 => x"00000000",
    25203 => x"00000000", 25204 => x"00000000", 25205 => x"00000000",
    25206 => x"00000000", 25207 => x"00000000", 25208 => x"00000000",
    25209 => x"00000000", 25210 => x"00000000", 25211 => x"00000000",
    25212 => x"00000000", 25213 => x"00000000", 25214 => x"00000000",
    25215 => x"00000000", 25216 => x"00000000", 25217 => x"00000000",
    25218 => x"00000000", 25219 => x"00000000", 25220 => x"00000000",
    25221 => x"00000000", 25222 => x"00000000", 25223 => x"00000000",
    25224 => x"00000000", 25225 => x"00000000", 25226 => x"00000000",
    25227 => x"00000000", 25228 => x"00000000", 25229 => x"00000000",
    25230 => x"00000000", 25231 => x"00000000", 25232 => x"00000000",
    25233 => x"00000000", 25234 => x"00000000", 25235 => x"00000000",
    25236 => x"00000000", 25237 => x"00000000", 25238 => x"00000000",
    25239 => x"00000000", 25240 => x"00000000", 25241 => x"00000000",
    25242 => x"00000000", 25243 => x"00000000", 25244 => x"00000000",
    25245 => x"00000000", 25246 => x"00000000", 25247 => x"00000000",
    25248 => x"00000000", 25249 => x"00000000", 25250 => x"00000000",
    25251 => x"00000000", 25252 => x"00000000", 25253 => x"00000000",
    25254 => x"00000000", 25255 => x"00000000", 25256 => x"00000000",
    25257 => x"00000000", 25258 => x"00000000", 25259 => x"00000000",
    25260 => x"00000000", 25261 => x"00000000", 25262 => x"00000000",
    25263 => x"00000000", 25264 => x"00000000", 25265 => x"00000000",
    25266 => x"00000000", 25267 => x"00000000", 25268 => x"00000000",
    25269 => x"00000000", 25270 => x"00000000", 25271 => x"00000000",
    25272 => x"00000000", 25273 => x"00000000", 25274 => x"00000000",
    25275 => x"00000000", 25276 => x"00000000", 25277 => x"00000000",
    25278 => x"00000000", 25279 => x"00000000", 25280 => x"00000000",
    25281 => x"00000000", 25282 => x"00000000", 25283 => x"00000000",
    25284 => x"00000000", 25285 => x"00000000", 25286 => x"00000000",
    25287 => x"00000000", 25288 => x"00000000", 25289 => x"00000000",
    25290 => x"00000000", 25291 => x"00000000", 25292 => x"00000000",
    25293 => x"00000000", 25294 => x"00000000", 25295 => x"00000000",
    25296 => x"00000000", 25297 => x"00000000", 25298 => x"00000000",
    25299 => x"00000000", 25300 => x"00000000", 25301 => x"00000000",
    25302 => x"00000000", 25303 => x"00000000", 25304 => x"00000000",
    25305 => x"00000000", 25306 => x"00000000", 25307 => x"00000000",
    25308 => x"00000000", 25309 => x"00000000", 25310 => x"00000000",
    25311 => x"00000000", 25312 => x"00000000", 25313 => x"00000000",
    25314 => x"00000000", 25315 => x"00000000", 25316 => x"00000000",
    25317 => x"00000000", 25318 => x"00000000", 25319 => x"00000000",
    25320 => x"00000000", 25321 => x"00000000", 25322 => x"00000000",
    25323 => x"00000000", 25324 => x"00000000", 25325 => x"00000000",
    25326 => x"00000000", 25327 => x"00000000", 25328 => x"00000000",
    25329 => x"00000000", 25330 => x"00000000", 25331 => x"00000000",
    25332 => x"00000000", 25333 => x"00000000", 25334 => x"00000000",
    25335 => x"00000000", 25336 => x"00000000", 25337 => x"00000000",
    25338 => x"00000000", 25339 => x"00000000", 25340 => x"00000000",
    25341 => x"00000000", 25342 => x"00000000", 25343 => x"00000000",
    25344 => x"00000000", 25345 => x"00000000", 25346 => x"00000000",
    25347 => x"00000000", 25348 => x"00000000", 25349 => x"00000000",
    25350 => x"00000000", 25351 => x"00000000", 25352 => x"00000000",
    25353 => x"00000000", 25354 => x"00000000", 25355 => x"00000000",
    25356 => x"00000000", 25357 => x"00000000", 25358 => x"00000000",
    25359 => x"00000000", 25360 => x"00000000", 25361 => x"00000000",
    25362 => x"00000000", 25363 => x"00000000", 25364 => x"00000000",
    25365 => x"00000000", 25366 => x"00000000", 25367 => x"00000000",
    25368 => x"00000000", 25369 => x"00000000", 25370 => x"00000000",
    25371 => x"00000000", 25372 => x"00000000", 25373 => x"00000000",
    25374 => x"00000000", 25375 => x"00000000", 25376 => x"00000000",
    25377 => x"00000000", 25378 => x"00000000", 25379 => x"00000000",
    25380 => x"00000000", 25381 => x"00000000", 25382 => x"00000000",
    25383 => x"00000000", 25384 => x"00000000", 25385 => x"00000000",
    25386 => x"00000000", 25387 => x"00000000", 25388 => x"00000000",
    25389 => x"00000000", 25390 => x"00000000", 25391 => x"00000000",
    25392 => x"00000000", 25393 => x"00000000", 25394 => x"00000000",
    25395 => x"00000000", 25396 => x"00000000", 25397 => x"00000000",
    25398 => x"00000000", 25399 => x"00000000", 25400 => x"00000000",
    25401 => x"00000000", 25402 => x"00000000", 25403 => x"00000000",
    25404 => x"00000000", 25405 => x"00000000", 25406 => x"00000000",
    25407 => x"00000000", 25408 => x"00000000", 25409 => x"00000000",
    25410 => x"00000000", 25411 => x"00000000", 25412 => x"00000000",
    25413 => x"00000000", 25414 => x"00000000", 25415 => x"00000000",
    25416 => x"00000000", 25417 => x"00000000", 25418 => x"00000000",
    25419 => x"00000000", 25420 => x"00000000", 25421 => x"00000000",
    25422 => x"00000000", 25423 => x"00000000", 25424 => x"00000000",
    25425 => x"00000000", 25426 => x"00000000", 25427 => x"00000000",
    25428 => x"00000000", 25429 => x"00000000", 25430 => x"00000000",
    25431 => x"00000000", 25432 => x"00000000", 25433 => x"00000000",
    25434 => x"00000000", 25435 => x"00000000", 25436 => x"00000000",
    25437 => x"00000000", 25438 => x"00000000", 25439 => x"00000000",
    25440 => x"00000000", 25441 => x"00000000", 25442 => x"00000000",
    25443 => x"00000000", 25444 => x"00000000", 25445 => x"00000000",
    25446 => x"00000000", 25447 => x"00000000", 25448 => x"00000000",
    25449 => x"00000000", 25450 => x"00000000", 25451 => x"00000000",
    25452 => x"00000000", 25453 => x"00000000", 25454 => x"00000000",
    25455 => x"00000000", 25456 => x"00000000", 25457 => x"00000000",
    25458 => x"00000000", 25459 => x"00000000", 25460 => x"00000000",
    25461 => x"00000000", 25462 => x"00000000", 25463 => x"00000000",
    25464 => x"00000000", 25465 => x"00000000", 25466 => x"00000000",
    25467 => x"00000000", 25468 => x"00000000", 25469 => x"00000000",
    25470 => x"00000000", 25471 => x"00000000", 25472 => x"00000000",
    25473 => x"00000000", 25474 => x"00000000", 25475 => x"00000000",
    25476 => x"00000000", 25477 => x"00000000", 25478 => x"00000000",
    25479 => x"00000000", 25480 => x"00000000", 25481 => x"00000000",
    25482 => x"00000000", 25483 => x"00000000", 25484 => x"00000000",
    25485 => x"00000000", 25486 => x"00000000", 25487 => x"00000000",
    25488 => x"00000000", 25489 => x"00000000", 25490 => x"00000000",
    25491 => x"00000000", 25492 => x"00000000", 25493 => x"00000000",
    25494 => x"00000000", 25495 => x"00000000", 25496 => x"00000000",
    25497 => x"00000000", 25498 => x"00000000", 25499 => x"00000000",
    25500 => x"00000000", 25501 => x"00000000", 25502 => x"00000000",
    25503 => x"00000000", 25504 => x"00000000", 25505 => x"00000000",
    25506 => x"00000000", 25507 => x"00000000", 25508 => x"00000000",
    25509 => x"00000000", 25510 => x"00000000", 25511 => x"00000000",
    25512 => x"00000000", 25513 => x"00000000", 25514 => x"00000000",
    25515 => x"00000000", 25516 => x"00000000", 25517 => x"00000000",
    25518 => x"00000000", 25519 => x"00000000", 25520 => x"00000000",
    25521 => x"00000000", 25522 => x"00000000", 25523 => x"00000000",
    25524 => x"00000000", 25525 => x"00000000", 25526 => x"00000000",
    25527 => x"00000000", 25528 => x"00000000", 25529 => x"00000000",
    25530 => x"00000000", 25531 => x"00000000", 25532 => x"00000000",
    25533 => x"00000000", 25534 => x"00000000", 25535 => x"00000000",
    25536 => x"00000000", 25537 => x"00000000", 25538 => x"00000000",
    25539 => x"00000000", 25540 => x"00000000", 25541 => x"00000000",
    25542 => x"00000000", 25543 => x"00000000", 25544 => x"00000000",
    25545 => x"00000000", 25546 => x"00000000", 25547 => x"00000000",
    25548 => x"00000000", 25549 => x"00000000", 25550 => x"00000000",
    25551 => x"00000000", 25552 => x"00000000", 25553 => x"00000000",
    25554 => x"00000000", 25555 => x"00000000", 25556 => x"00000000",
    25557 => x"00000000", 25558 => x"00000000", 25559 => x"00000000",
    25560 => x"00000000", 25561 => x"00000000", 25562 => x"00000000",
    25563 => x"00000000", 25564 => x"00000000", 25565 => x"00000000",
    25566 => x"00000000", 25567 => x"00000000", 25568 => x"00000000",
    25569 => x"00000000", 25570 => x"00000000", 25571 => x"00000000",
    25572 => x"00000000", 25573 => x"00000000", 25574 => x"00000000",
    25575 => x"00000000", 25576 => x"00000000", 25577 => x"00000000",
    25578 => x"00000000", 25579 => x"00000000", 25580 => x"00000000",
    25581 => x"00000000", 25582 => x"00000000", 25583 => x"00000000",
    25584 => x"00000000", 25585 => x"00000000", 25586 => x"00000000",
    25587 => x"00000000", 25588 => x"00000000", 25589 => x"00000000",
    25590 => x"00000000", 25591 => x"00000000", 25592 => x"00000000",
    25593 => x"00000000", 25594 => x"00000000", 25595 => x"00000000",
    25596 => x"00000000", 25597 => x"00000000", 25598 => x"00000000",
    25599 => x"00000000", 25600 => x"00000000", 25601 => x"00000000",
    25602 => x"00000000", 25603 => x"00000000", 25604 => x"00000000",
    25605 => x"00000000", 25606 => x"00000000", 25607 => x"00000000",
    25608 => x"00000000", 25609 => x"00000000", 25610 => x"00000000",
    25611 => x"00000000", 25612 => x"00000000", 25613 => x"00000000",
    25614 => x"00000000", 25615 => x"00000000", 25616 => x"00000000",
    25617 => x"00000000", 25618 => x"00000000", 25619 => x"00000000",
    25620 => x"00000000", 25621 => x"00000000", 25622 => x"00000000",
    25623 => x"00000000", 25624 => x"00000000", 25625 => x"00000000",
    25626 => x"00000000", 25627 => x"00000000", 25628 => x"00000000",
    25629 => x"00000000", 25630 => x"00000000", 25631 => x"00000000",
    25632 => x"00000000", 25633 => x"00000000", 25634 => x"00000000",
    25635 => x"00000000", 25636 => x"00000000", 25637 => x"00000000",
    25638 => x"00000000", 25639 => x"00000000", 25640 => x"00000000",
    25641 => x"00000000", 25642 => x"00000000", 25643 => x"00000000",
    25644 => x"00000000", 25645 => x"00000000", 25646 => x"00000000",
    25647 => x"00000000", 25648 => x"00000000", 25649 => x"00000000",
    25650 => x"00000000", 25651 => x"00000000", 25652 => x"00000000",
    25653 => x"00000000", 25654 => x"00000000", 25655 => x"00000000",
    25656 => x"00000000", 25657 => x"00000000", 25658 => x"00000000",
    25659 => x"00000000", 25660 => x"00000000", 25661 => x"00000000",
    25662 => x"00000000", 25663 => x"00000000", 25664 => x"00000000",
    25665 => x"00000000", 25666 => x"00000000", 25667 => x"00000000",
    25668 => x"00000000", 25669 => x"00000000", 25670 => x"00000000",
    25671 => x"00000000", 25672 => x"00000000", 25673 => x"00000000",
    25674 => x"00000000", 25675 => x"00000000", 25676 => x"00000000",
    25677 => x"00000000", 25678 => x"00000000", 25679 => x"00000000",
    25680 => x"00000000", 25681 => x"00000000", 25682 => x"00000000",
    25683 => x"00000000", 25684 => x"00000000", 25685 => x"00000000",
    25686 => x"00000000", 25687 => x"00000000", 25688 => x"00000000",
    25689 => x"00000000", 25690 => x"00000000", 25691 => x"00000000",
    25692 => x"00000000", 25693 => x"00000000", 25694 => x"00000000",
    25695 => x"00000000", 25696 => x"00000000", 25697 => x"00000000",
    25698 => x"00000000", 25699 => x"00000000", 25700 => x"00000000",
    25701 => x"00000000", 25702 => x"00000000", 25703 => x"00000000",
    25704 => x"00000000", 25705 => x"00000000", 25706 => x"00000000",
    25707 => x"00000000", 25708 => x"00000000", 25709 => x"00000000",
    25710 => x"00000000", 25711 => x"00000000", 25712 => x"00000000",
    25713 => x"00000000", 25714 => x"00000000", 25715 => x"00000000",
    25716 => x"00000000", 25717 => x"00000000", 25718 => x"00000000",
    25719 => x"00000000", 25720 => x"00000000", 25721 => x"00000000",
    25722 => x"00000000", 25723 => x"00000000", 25724 => x"00000000",
    25725 => x"00000000", 25726 => x"00000000", 25727 => x"00000000",
    25728 => x"00000000", 25729 => x"00000000", 25730 => x"00000000",
    25731 => x"00000000", 25732 => x"00000000", 25733 => x"00000000",
    25734 => x"00000000", 25735 => x"00000000", 25736 => x"00000000",
    25737 => x"00000000", 25738 => x"00000000", 25739 => x"00000000",
    25740 => x"00000000", 25741 => x"00000000", 25742 => x"00000000",
    25743 => x"00000000", 25744 => x"00000000", 25745 => x"00000000",
    25746 => x"00000000", 25747 => x"00000000", 25748 => x"00000000",
    25749 => x"00000000", 25750 => x"00000000", 25751 => x"00000000",
    25752 => x"00000000", 25753 => x"00000000", 25754 => x"00000000",
    25755 => x"00000000", 25756 => x"00000000", 25757 => x"00000000",
    25758 => x"00000000", 25759 => x"00000000", 25760 => x"00000000",
    25761 => x"00000000", 25762 => x"00000000", 25763 => x"00000000",
    25764 => x"00000000", 25765 => x"00000000", 25766 => x"00000000",
    25767 => x"00000000", 25768 => x"00000000", 25769 => x"00000000",
    25770 => x"00000000", 25771 => x"00000000", 25772 => x"00000000",
    25773 => x"00000000", 25774 => x"00000000", 25775 => x"00000000",
    25776 => x"00000000", 25777 => x"00000000", 25778 => x"00000000",
    25779 => x"00000000", 25780 => x"00000000", 25781 => x"00000000",
    25782 => x"00000000", 25783 => x"00000000", 25784 => x"00000000",
    25785 => x"00000000", 25786 => x"00000000", 25787 => x"00000000",
    25788 => x"00000000", 25789 => x"00000000", 25790 => x"00000000",
    25791 => x"00000000", 25792 => x"00000000", 25793 => x"00000000",
    25794 => x"00000000", 25795 => x"00000000", 25796 => x"00000000",
    25797 => x"00000000", 25798 => x"00000000", 25799 => x"00000000",
    25800 => x"00000000", 25801 => x"00000000", 25802 => x"00000000",
    25803 => x"00000000", 25804 => x"00000000", 25805 => x"00000000",
    25806 => x"00000000", 25807 => x"00000000", 25808 => x"00000000",
    25809 => x"00000000", 25810 => x"00000000", 25811 => x"00000000",
    25812 => x"00000000", 25813 => x"00000000", 25814 => x"00000000",
    25815 => x"00000000", 25816 => x"00000000", 25817 => x"00000000",
    25818 => x"00000000", 25819 => x"00000000", 25820 => x"00000000",
    25821 => x"00000000", 25822 => x"00000000", 25823 => x"00000000",
    25824 => x"00000000", 25825 => x"00000000", 25826 => x"00000000",
    25827 => x"00000000", 25828 => x"00000000", 25829 => x"00000000",
    25830 => x"00000000", 25831 => x"00000000", 25832 => x"00000000",
    25833 => x"00000000", 25834 => x"00000000", 25835 => x"00000000",
    25836 => x"00000000", 25837 => x"00000000", 25838 => x"00000000",
    25839 => x"00000000", 25840 => x"00000000", 25841 => x"00000000",
    25842 => x"00000000", 25843 => x"00000000", 25844 => x"00000000",
    25845 => x"00000000", 25846 => x"00000000", 25847 => x"00000000",
    25848 => x"00000000", 25849 => x"00000000", 25850 => x"00000000",
    25851 => x"00000000", 25852 => x"00000000", 25853 => x"00000000",
    25854 => x"00000000", 25855 => x"00000000", 25856 => x"00000000",
    25857 => x"00000000", 25858 => x"00000000", 25859 => x"00000000",
    25860 => x"00000000", 25861 => x"00000000", 25862 => x"00000000",
    25863 => x"00000000", 25864 => x"00000000", 25865 => x"00000000",
    25866 => x"00000000", 25867 => x"00000000", 25868 => x"00000000",
    25869 => x"00000000", 25870 => x"00000000", 25871 => x"00000000",
    25872 => x"00000000", 25873 => x"00000000", 25874 => x"00000000",
    25875 => x"00000000", 25876 => x"00000000", 25877 => x"00000000",
    25878 => x"00000000", 25879 => x"00000000", 25880 => x"00000000",
    25881 => x"00000000", 25882 => x"00000000", 25883 => x"00000000",
    25884 => x"00000000", 25885 => x"00000000", 25886 => x"00000000",
    25887 => x"00000000", 25888 => x"00000000", 25889 => x"00000000",
    25890 => x"00000000", 25891 => x"00000000", 25892 => x"00000000",
    25893 => x"00000000", 25894 => x"00000000", 25895 => x"00000000",
    25896 => x"00000000", 25897 => x"00000000", 25898 => x"00000000",
    25899 => x"00000000", 25900 => x"00000000", 25901 => x"00000000",
    25902 => x"00000000", 25903 => x"00000000", 25904 => x"00000000",
    25905 => x"00000000", 25906 => x"00000000", 25907 => x"00000000",
    25908 => x"00000000", 25909 => x"00000000", 25910 => x"00000000",
    25911 => x"00000000", 25912 => x"00000000", 25913 => x"00000000",
    25914 => x"00000000", 25915 => x"00000000", 25916 => x"00000000",
    25917 => x"00000000", 25918 => x"00000000", 25919 => x"00000000",
    25920 => x"00000000", 25921 => x"00000000", 25922 => x"00000000",
    25923 => x"00000000", 25924 => x"00000000", 25925 => x"00000000",
    25926 => x"00000000", 25927 => x"00000000", 25928 => x"00000000",
    25929 => x"00000000", 25930 => x"00000000", 25931 => x"00000000",
    25932 => x"00000000", 25933 => x"00000000", 25934 => x"00000000",
    25935 => x"00000000", 25936 => x"00000000", 25937 => x"00000000",
    25938 => x"00000000", 25939 => x"00000000", 25940 => x"00000000",
    25941 => x"00000000", 25942 => x"00000000", 25943 => x"00000000",
    25944 => x"00000000", 25945 => x"00000000", 25946 => x"00000000",
    25947 => x"00000000", 25948 => x"00000000", 25949 => x"00000000",
    25950 => x"00000000", 25951 => x"00000000", 25952 => x"00000000",
    25953 => x"00000000", 25954 => x"00000000", 25955 => x"00000000",
    25956 => x"00000000", 25957 => x"00000000", 25958 => x"00000000",
    25959 => x"00000000", 25960 => x"00000000", 25961 => x"00000000",
    25962 => x"00000000", 25963 => x"00000000", 25964 => x"00000000",
    25965 => x"00000000", 25966 => x"00000000", 25967 => x"00000000",
    25968 => x"00000000", 25969 => x"00000000", 25970 => x"00000000",
    25971 => x"00000000", 25972 => x"00000000", 25973 => x"00000000",
    25974 => x"00000000", 25975 => x"00000000", 25976 => x"00000000",
    25977 => x"00000000", 25978 => x"00000000", 25979 => x"00000000",
    25980 => x"00000000", 25981 => x"00000000", 25982 => x"00000000",
    25983 => x"00000000", 25984 => x"00000000", 25985 => x"00000000",
    25986 => x"00000000", 25987 => x"00000000", 25988 => x"00000000",
    25989 => x"00000000", 25990 => x"00000000", 25991 => x"00000000",
    25992 => x"00000000", 25993 => x"00000000", 25994 => x"00000000",
    25995 => x"00000000", 25996 => x"00000000", 25997 => x"00000000",
    25998 => x"00000000", 25999 => x"00000000", 26000 => x"00000000",
    26001 => x"00000000", 26002 => x"00000000", 26003 => x"00000000",
    26004 => x"00000000", 26005 => x"00000000", 26006 => x"00000000",
    26007 => x"00000000", 26008 => x"00000000", 26009 => x"00000000",
    26010 => x"00000000", 26011 => x"00000000", 26012 => x"00000000",
    26013 => x"00000000", 26014 => x"00000000", 26015 => x"00000000",
    26016 => x"00000000", 26017 => x"00000000", 26018 => x"00000000",
    26019 => x"00000000", 26020 => x"00000000", 26021 => x"00000000",
    26022 => x"00000000", 26023 => x"00000000", 26024 => x"00000000",
    26025 => x"00000000", 26026 => x"00000000", 26027 => x"00000000",
    26028 => x"00000000", 26029 => x"00000000", 26030 => x"00000000",
    26031 => x"00000000", 26032 => x"00000000", 26033 => x"00000000",
    26034 => x"00000000", 26035 => x"00000000", 26036 => x"00000000",
    26037 => x"00000000", 26038 => x"00000000", 26039 => x"00000000",
    26040 => x"00000000", 26041 => x"00000000", 26042 => x"00000000",
    26043 => x"00000000", 26044 => x"00000000", 26045 => x"00000000",
    26046 => x"00000000", 26047 => x"00000000", 26048 => x"00000000",
    26049 => x"00000000", 26050 => x"00000000", 26051 => x"00000000",
    26052 => x"00000000", 26053 => x"00000000", 26054 => x"00000000",
    26055 => x"00000000", 26056 => x"00000000", 26057 => x"00000000",
    26058 => x"00000000", 26059 => x"00000000", 26060 => x"00000000",
    26061 => x"00000000", 26062 => x"00000000", 26063 => x"00000000",
    26064 => x"00000000", 26065 => x"00000000", 26066 => x"00000000",
    26067 => x"00000000", 26068 => x"00000000", 26069 => x"00000000",
    26070 => x"00000000", 26071 => x"00000000", 26072 => x"00000000",
    26073 => x"00000000", 26074 => x"00000000", 26075 => x"00000000",
    26076 => x"00000000", 26077 => x"00000000", 26078 => x"00000000",
    26079 => x"00000000", 26080 => x"00000000", 26081 => x"00000000",
    26082 => x"00000000", 26083 => x"00000000", 26084 => x"00000000",
    26085 => x"00000000", 26086 => x"00000000", 26087 => x"00000000",
    26088 => x"00000000", 26089 => x"00000000", 26090 => x"00000000",
    26091 => x"00000000", 26092 => x"00000000", 26093 => x"00000000",
    26094 => x"00000000", 26095 => x"00000000", 26096 => x"00000000",
    26097 => x"00000000", 26098 => x"00000000", 26099 => x"00000000",
    26100 => x"00000000", 26101 => x"00000000", 26102 => x"00000000",
    26103 => x"00000000", 26104 => x"00000000", 26105 => x"00000000",
    26106 => x"00000000", 26107 => x"00000000", 26108 => x"00000000",
    26109 => x"00000000", 26110 => x"00000000", 26111 => x"00000000",
    26112 => x"00000000", 26113 => x"00000000", 26114 => x"00000000",
    26115 => x"00000000", 26116 => x"00000000", 26117 => x"00000000",
    26118 => x"00000000", 26119 => x"00000000", 26120 => x"00000000",
    26121 => x"00000000", 26122 => x"00000000", 26123 => x"00000000",
    26124 => x"00000000", 26125 => x"00000000", 26126 => x"00000000",
    26127 => x"00000000", 26128 => x"00000000", 26129 => x"00000000",
    26130 => x"00000000", 26131 => x"00000000", 26132 => x"00000000",
    26133 => x"00000000", 26134 => x"00000000", 26135 => x"00000000",
    26136 => x"00000000", 26137 => x"00000000", 26138 => x"00000000",
    26139 => x"00000000", 26140 => x"00000000", 26141 => x"00000000",
    26142 => x"00000000", 26143 => x"00000000", 26144 => x"00000000",
    26145 => x"00000000", 26146 => x"00000000", 26147 => x"00000000",
    26148 => x"00000000", 26149 => x"00000000", 26150 => x"00000000",
    26151 => x"00000000", 26152 => x"00000000", 26153 => x"00000000",
    26154 => x"00000000", 26155 => x"00000000", 26156 => x"00000000",
    26157 => x"00000000", 26158 => x"00000000", 26159 => x"00000000",
    26160 => x"00000000", 26161 => x"00000000", 26162 => x"00000000",
    26163 => x"00000000", 26164 => x"00000000", 26165 => x"00000000",
    26166 => x"00000000", 26167 => x"00000000", 26168 => x"00000000",
    26169 => x"00000000", 26170 => x"00000000", 26171 => x"00000000",
    26172 => x"00000000", 26173 => x"00000000", 26174 => x"00000000",
    26175 => x"00000000", 26176 => x"00000000", 26177 => x"00000000",
    26178 => x"00000000", 26179 => x"00000000", 26180 => x"00000000",
    26181 => x"00000000", 26182 => x"00000000", 26183 => x"00000000",
    26184 => x"00000000", 26185 => x"00000000", 26186 => x"00000000",
    26187 => x"00000000", 26188 => x"00000000", 26189 => x"00000000",
    26190 => x"00000000", 26191 => x"00000000", 26192 => x"00000000",
    26193 => x"00000000", 26194 => x"00000000", 26195 => x"00000000",
    26196 => x"00000000", 26197 => x"00000000", 26198 => x"00000000",
    26199 => x"00000000", 26200 => x"00000000", 26201 => x"00000000",
    26202 => x"00000000", 26203 => x"00000000", 26204 => x"00000000",
    26205 => x"00000000", 26206 => x"00000000", 26207 => x"00000000",
    26208 => x"00000000", 26209 => x"00000000", 26210 => x"00000000",
    26211 => x"00000000", 26212 => x"00000000", 26213 => x"00000000",
    26214 => x"00000000", 26215 => x"00000000", 26216 => x"00000000",
    26217 => x"00000000", 26218 => x"00000000", 26219 => x"00000000",
    26220 => x"00000000", 26221 => x"00000000", 26222 => x"00000000",
    26223 => x"00000000", 26224 => x"00000000", 26225 => x"00000000",
    26226 => x"00000000", 26227 => x"00000000", 26228 => x"00000000",
    26229 => x"00000000", 26230 => x"00000000", 26231 => x"00000000",
    26232 => x"00000000", 26233 => x"00000000", 26234 => x"00000000",
    26235 => x"00000000", 26236 => x"00000000", 26237 => x"00000000",
    26238 => x"00000000", 26239 => x"00000000", 26240 => x"00000000",
    26241 => x"00000000", 26242 => x"00000000", 26243 => x"00000000",
    26244 => x"00000000", 26245 => x"00000000", 26246 => x"00000000",
    26247 => x"00000000", 26248 => x"00000000", 26249 => x"00000000",
    26250 => x"00000000", 26251 => x"00000000", 26252 => x"00000000",
    26253 => x"00000000", 26254 => x"00000000", 26255 => x"00000000",
    26256 => x"00000000", 26257 => x"00000000", 26258 => x"00000000",
    26259 => x"00000000", 26260 => x"00000000", 26261 => x"00000000",
    26262 => x"00000000", 26263 => x"00000000", 26264 => x"00000000",
    26265 => x"00000000", 26266 => x"00000000", 26267 => x"00000000",
    26268 => x"00000000", 26269 => x"00000000", 26270 => x"00000000",
    26271 => x"00000000", 26272 => x"00000000", 26273 => x"00000000",
    26274 => x"00000000", 26275 => x"00000000", 26276 => x"00000000",
    26277 => x"00000000", 26278 => x"00000000", 26279 => x"00000000",
    26280 => x"00000000", 26281 => x"00000000", 26282 => x"00000000",
    26283 => x"00000000", 26284 => x"00000000", 26285 => x"00000000",
    26286 => x"00000000", 26287 => x"00000000", 26288 => x"00000000",
    26289 => x"00000000", 26290 => x"00000000", 26291 => x"00000000",
    26292 => x"00000000", 26293 => x"00000000", 26294 => x"00000000",
    26295 => x"00000000", 26296 => x"00000000", 26297 => x"00000000",
    26298 => x"00000000", 26299 => x"00000000", 26300 => x"00000000",
    26301 => x"00000000", 26302 => x"00000000", 26303 => x"00000000",
    26304 => x"00000000", 26305 => x"00000000", 26306 => x"00000000",
    26307 => x"00000000", 26308 => x"00000000", 26309 => x"00000000",
    26310 => x"00000000", 26311 => x"00000000", 26312 => x"00000000",
    26313 => x"00000000", 26314 => x"00000000", 26315 => x"00000000",
    26316 => x"00000000", 26317 => x"00000000", 26318 => x"00000000",
    26319 => x"00000000", 26320 => x"00000000", 26321 => x"00000000",
    26322 => x"00000000", 26323 => x"00000000", 26324 => x"00000000",
    26325 => x"00000000", 26326 => x"00000000", 26327 => x"00000000",
    26328 => x"00000000", 26329 => x"00000000", 26330 => x"00000000",
    26331 => x"00000000", 26332 => x"00000000", 26333 => x"00000000",
    26334 => x"00000000", 26335 => x"00000000", 26336 => x"00000000",
    26337 => x"00000000", 26338 => x"00000000", 26339 => x"00000000",
    26340 => x"00000000", 26341 => x"00000000", 26342 => x"00000000",
    26343 => x"00000000", 26344 => x"00000000", 26345 => x"00000000",
    26346 => x"00000000", 26347 => x"00000000", 26348 => x"00000000",
    26349 => x"00000000", 26350 => x"00000000", 26351 => x"00000000",
    26352 => x"00000000", 26353 => x"00000000", 26354 => x"00000000",
    26355 => x"00000000", 26356 => x"00000000", 26357 => x"00000000",
    26358 => x"00000000", 26359 => x"00000000", 26360 => x"00000000",
    26361 => x"00000000", 26362 => x"00000000", 26363 => x"00000000",
    26364 => x"00000000", 26365 => x"00000000", 26366 => x"00000000",
    26367 => x"00000000", 26368 => x"00000000", 26369 => x"00000000",
    26370 => x"00000000", 26371 => x"00000000", 26372 => x"00000000",
    26373 => x"00000000", 26374 => x"00000000", 26375 => x"00000000",
    26376 => x"00000000", 26377 => x"00000000", 26378 => x"00000000",
    26379 => x"00000000", 26380 => x"00000000", 26381 => x"00000000",
    26382 => x"00000000", 26383 => x"00000000", 26384 => x"00000000",
    26385 => x"00000000", 26386 => x"00000000", 26387 => x"00000000",
    26388 => x"00000000", 26389 => x"00000000", 26390 => x"00000000",
    26391 => x"00000000", 26392 => x"00000000", 26393 => x"00000000",
    26394 => x"00000000", 26395 => x"00000000", 26396 => x"00000000",
    26397 => x"00000000", 26398 => x"00000000", 26399 => x"00000000",
    26400 => x"00000000", 26401 => x"00000000", 26402 => x"00000000",
    26403 => x"00000000", 26404 => x"00000000", 26405 => x"00000000",
    26406 => x"00000000", 26407 => x"00000000", 26408 => x"00000000",
    26409 => x"00000000", 26410 => x"00000000", 26411 => x"00000000",
    26412 => x"00000000", 26413 => x"00000000", 26414 => x"00000000",
    26415 => x"00000000", 26416 => x"00000000", 26417 => x"00000000",
    26418 => x"00000000", 26419 => x"00000000", 26420 => x"00000000",
    26421 => x"00000000", 26422 => x"00000000", 26423 => x"00000000",
    26424 => x"00000000", 26425 => x"00000000", 26426 => x"00000000",
    26427 => x"00000000", 26428 => x"00000000", 26429 => x"00000000",
    26430 => x"00000000", 26431 => x"00000000", 26432 => x"00000000",
    26433 => x"00000000", 26434 => x"00000000", 26435 => x"00000000",
    26436 => x"00000000", 26437 => x"00000000", 26438 => x"00000000",
    26439 => x"00000000", 26440 => x"00000000", 26441 => x"00000000",
    26442 => x"00000000", 26443 => x"00000000", 26444 => x"00000000",
    26445 => x"00000000", 26446 => x"00000000", 26447 => x"00000000",
    26448 => x"00000000", 26449 => x"00000000", 26450 => x"00000000",
    26451 => x"00000000", 26452 => x"00000000", 26453 => x"00000000",
    26454 => x"00000000", 26455 => x"00000000", 26456 => x"00000000",
    26457 => x"00000000", 26458 => x"00000000", 26459 => x"00000000",
    26460 => x"00000000", 26461 => x"00000000", 26462 => x"00000000",
    26463 => x"00000000", 26464 => x"00000000", 26465 => x"00000000",
    26466 => x"00000000", 26467 => x"00000000", 26468 => x"00000000",
    26469 => x"00000000", 26470 => x"00000000", 26471 => x"00000000",
    26472 => x"00000000", 26473 => x"00000000", 26474 => x"00000000",
    26475 => x"00000000", 26476 => x"00000000", 26477 => x"00000000",
    26478 => x"00000000", 26479 => x"00000000", 26480 => x"00000000",
    26481 => x"00000000", 26482 => x"00000000", 26483 => x"00000000",
    26484 => x"00000000", 26485 => x"00000000", 26486 => x"00000000",
    26487 => x"00000000", 26488 => x"00000000", 26489 => x"00000000",
    26490 => x"00000000", 26491 => x"00000000", 26492 => x"00000000",
    26493 => x"00000000", 26494 => x"00000000", 26495 => x"00000000",
    26496 => x"00000000", 26497 => x"00000000", 26498 => x"00000000",
    26499 => x"00000000", 26500 => x"00000000", 26501 => x"00000000",
    26502 => x"00000000", 26503 => x"00000000", 26504 => x"00000000",
    26505 => x"00000000", 26506 => x"00000000", 26507 => x"00000000",
    26508 => x"00000000", 26509 => x"00000000", 26510 => x"00000000",
    26511 => x"00000000", 26512 => x"00000000", 26513 => x"00000000",
    26514 => x"00000000", 26515 => x"00000000", 26516 => x"00000000",
    26517 => x"00000000", 26518 => x"00000000", 26519 => x"00000000",
    26520 => x"00000000", 26521 => x"00000000", 26522 => x"00000000",
    26523 => x"00000000", 26524 => x"00000000", 26525 => x"00000000",
    26526 => x"00000000", 26527 => x"00000000", 26528 => x"00000000",
    26529 => x"00000000", 26530 => x"00000000", 26531 => x"00000000",
    26532 => x"00000000", 26533 => x"00000000", 26534 => x"00000000",
    26535 => x"00000000", 26536 => x"00000000", 26537 => x"00000000",
    26538 => x"00000000", 26539 => x"00000000", 26540 => x"00000000",
    26541 => x"00000000", 26542 => x"00000000", 26543 => x"00000000",
    26544 => x"00000000", 26545 => x"00000000", 26546 => x"00000000",
    26547 => x"00000000", 26548 => x"00000000", 26549 => x"00000000",
    26550 => x"00000000", 26551 => x"00000000", 26552 => x"00000000",
    26553 => x"00000000", 26554 => x"00000000", 26555 => x"00000000",
    26556 => x"00000000", 26557 => x"00000000", 26558 => x"00000000",
    26559 => x"00000000", 26560 => x"00000000", 26561 => x"00000000",
    26562 => x"00000000", 26563 => x"00000000", 26564 => x"00000000",
    26565 => x"00000000", 26566 => x"00000000", 26567 => x"00000000",
    26568 => x"00000000", 26569 => x"00000000", 26570 => x"00000000",
    26571 => x"00000000", 26572 => x"00000000", 26573 => x"00000000",
    26574 => x"00000000", 26575 => x"00000000", 26576 => x"00000000",
    26577 => x"00000000", 26578 => x"00000000", 26579 => x"00000000",
    26580 => x"00000000", 26581 => x"00000000", 26582 => x"00000000",
    26583 => x"00000000", 26584 => x"00000000", 26585 => x"00000000",
    26586 => x"00000000", 26587 => x"00000000", 26588 => x"00000000",
    26589 => x"00000000", 26590 => x"00000000", 26591 => x"00000000",
    26592 => x"00000000", 26593 => x"00000000", 26594 => x"00000000",
    26595 => x"00000000", 26596 => x"00000000", 26597 => x"00000000",
    26598 => x"00000000", 26599 => x"00000000", 26600 => x"00000000",
    26601 => x"00000000", 26602 => x"00000000", 26603 => x"00000000",
    26604 => x"00000000", 26605 => x"00000000", 26606 => x"00000000",
    26607 => x"00000000", 26608 => x"00000000", 26609 => x"00000000",
    26610 => x"00000000", 26611 => x"00000000", 26612 => x"00000000",
    26613 => x"00000000", 26614 => x"00000000", 26615 => x"00000000",
    26616 => x"00000000", 26617 => x"00000000", 26618 => x"00000000",
    26619 => x"00000000", 26620 => x"00000000", 26621 => x"00000000",
    26622 => x"00000000", 26623 => x"00000000", 26624 => x"00000000",
    26625 => x"00000000", 26626 => x"00000000", 26627 => x"00000000",
    26628 => x"00000000", 26629 => x"00000000", 26630 => x"00000000",
    26631 => x"00000000", 26632 => x"00000000", 26633 => x"00000000",
    26634 => x"00000000", 26635 => x"00000000", 26636 => x"00000000",
    26637 => x"00000000", 26638 => x"00000000", 26639 => x"00000000",
    26640 => x"00000000", 26641 => x"00000000", 26642 => x"00000000",
    26643 => x"00000000", 26644 => x"00000000", 26645 => x"00000000",
    26646 => x"00000000", 26647 => x"00000000", 26648 => x"00000000",
    26649 => x"00000000", 26650 => x"00000000", 26651 => x"00000000",
    26652 => x"00000000", 26653 => x"00000000", 26654 => x"00000000",
    26655 => x"00000000", 26656 => x"00000000", 26657 => x"00000000",
    26658 => x"00000000", 26659 => x"00000000", 26660 => x"00000000",
    26661 => x"00000000", 26662 => x"00000000", 26663 => x"00000000",
    26664 => x"00000000", 26665 => x"00000000", 26666 => x"00000000",
    26667 => x"00000000", 26668 => x"00000000", 26669 => x"00000000",
    26670 => x"00000000", 26671 => x"00000000", 26672 => x"00000000",
    26673 => x"00000000", 26674 => x"00000000", 26675 => x"00000000",
    26676 => x"00000000", 26677 => x"00000000", 26678 => x"00000000",
    26679 => x"00000000", 26680 => x"00000000", 26681 => x"00000000",
    26682 => x"00000000", 26683 => x"00000000", 26684 => x"00000000",
    26685 => x"00000000", 26686 => x"00000000", 26687 => x"00000000",
    26688 => x"00000000", 26689 => x"00000000", 26690 => x"00000000",
    26691 => x"00000000", 26692 => x"00000000", 26693 => x"00000000",
    26694 => x"00000000", 26695 => x"00000000", 26696 => x"00000000",
    26697 => x"00000000", 26698 => x"00000000", 26699 => x"00000000",
    26700 => x"00000000", 26701 => x"00000000", 26702 => x"00000000",
    26703 => x"00000000", 26704 => x"00000000", 26705 => x"00000000",
    26706 => x"00000000", 26707 => x"00000000", 26708 => x"00000000",
    26709 => x"00000000", 26710 => x"00000000", 26711 => x"00000000",
    26712 => x"00000000", 26713 => x"00000000", 26714 => x"00000000",
    26715 => x"00000000", 26716 => x"00000000", 26717 => x"00000000",
    26718 => x"00000000", 26719 => x"00000000", 26720 => x"00000000",
    26721 => x"00000000", 26722 => x"00000000", 26723 => x"00000000",
    26724 => x"00000000", 26725 => x"00000000", 26726 => x"00000000",
    26727 => x"00000000", 26728 => x"00000000", 26729 => x"00000000",
    26730 => x"00000000", 26731 => x"00000000", 26732 => x"00000000",
    26733 => x"00000000", 26734 => x"00000000", 26735 => x"00000000",
    26736 => x"00000000", 26737 => x"00000000", 26738 => x"00000000",
    26739 => x"00000000", 26740 => x"00000000", 26741 => x"00000000",
    26742 => x"00000000", 26743 => x"00000000", 26744 => x"00000000",
    26745 => x"00000000", 26746 => x"00000000", 26747 => x"00000000",
    26748 => x"00000000", 26749 => x"00000000", 26750 => x"00000000",
    26751 => x"00000000", 26752 => x"00000000", 26753 => x"00000000",
    26754 => x"00000000", 26755 => x"00000000", 26756 => x"00000000",
    26757 => x"00000000", 26758 => x"00000000", 26759 => x"00000000",
    26760 => x"00000000", 26761 => x"00000000", 26762 => x"00000000",
    26763 => x"00000000", 26764 => x"00000000", 26765 => x"00000000",
    26766 => x"00000000", 26767 => x"00000000", 26768 => x"00000000",
    26769 => x"00000000", 26770 => x"00000000", 26771 => x"00000000",
    26772 => x"00000000", 26773 => x"00000000", 26774 => x"00000000",
    26775 => x"00000000", 26776 => x"00000000", 26777 => x"00000000",
    26778 => x"00000000", 26779 => x"00000000", 26780 => x"00000000",
    26781 => x"00000000", 26782 => x"00000000", 26783 => x"00000000",
    26784 => x"00000000", 26785 => x"00000000", 26786 => x"00000000",
    26787 => x"00000000", 26788 => x"00000000", 26789 => x"00000000",
    26790 => x"00000000", 26791 => x"00000000", 26792 => x"00000000",
    26793 => x"00000000", 26794 => x"00000000", 26795 => x"00000000",
    26796 => x"00000000", 26797 => x"00000000", 26798 => x"00000000",
    26799 => x"00000000", 26800 => x"00000000", 26801 => x"00000000",
    26802 => x"00000000", 26803 => x"00000000", 26804 => x"00000000",
    26805 => x"00000000", 26806 => x"00000000", 26807 => x"00000000",
    26808 => x"00000000", 26809 => x"00000000", 26810 => x"00000000",
    26811 => x"00000000", 26812 => x"00000000", 26813 => x"00000000",
    26814 => x"00000000", 26815 => x"00000000", 26816 => x"00000000",
    26817 => x"00000000", 26818 => x"00000000", 26819 => x"00000000",
    26820 => x"00000000", 26821 => x"00000000", 26822 => x"00000000",
    26823 => x"00000000", 26824 => x"00000000", 26825 => x"00000000",
    26826 => x"00000000", 26827 => x"00000000", 26828 => x"00000000",
    26829 => x"00000000", 26830 => x"00000000", 26831 => x"00000000",
    26832 => x"00000000", 26833 => x"00000000", 26834 => x"00000000",
    26835 => x"00000000", 26836 => x"00000000", 26837 => x"00000000",
    26838 => x"00000000", 26839 => x"00000000", 26840 => x"00000000",
    26841 => x"00000000", 26842 => x"00000000", 26843 => x"00000000",
    26844 => x"00000000", 26845 => x"00000000", 26846 => x"00000000",
    26847 => x"00000000", 26848 => x"00000000", 26849 => x"00000000",
    26850 => x"00000000", 26851 => x"00000000", 26852 => x"00000000",
    26853 => x"00000000", 26854 => x"00000000", 26855 => x"00000000",
    26856 => x"00000000", 26857 => x"00000000", 26858 => x"00000000",
    26859 => x"00000000", 26860 => x"00000000", 26861 => x"00000000",
    26862 => x"00000000", 26863 => x"00000000", 26864 => x"00000000",
    26865 => x"00000000", 26866 => x"00000000", 26867 => x"00000000",
    26868 => x"00000000", 26869 => x"00000000", 26870 => x"00000000",
    26871 => x"00000000", 26872 => x"00000000", 26873 => x"00000000",
    26874 => x"00000000", 26875 => x"00000000", 26876 => x"00000000",
    26877 => x"00000000", 26878 => x"00000000", 26879 => x"00000000",
    26880 => x"00000000", 26881 => x"00000000", 26882 => x"00000000",
    26883 => x"00000000", 26884 => x"00000000", 26885 => x"00000000",
    26886 => x"00000000", 26887 => x"00000000", 26888 => x"00000000",
    26889 => x"00000000", 26890 => x"00000000", 26891 => x"00000000",
    26892 => x"00000000", 26893 => x"00000000", 26894 => x"00000000",
    26895 => x"00000000", 26896 => x"00000000", 26897 => x"00000000",
    26898 => x"00000000", 26899 => x"00000000", 26900 => x"00000000",
    26901 => x"00000000", 26902 => x"00000000", 26903 => x"00000000",
    26904 => x"00000000", 26905 => x"00000000", 26906 => x"00000000",
    26907 => x"00000000", 26908 => x"00000000", 26909 => x"00000000",
    26910 => x"00000000", 26911 => x"00000000", 26912 => x"00000000",
    26913 => x"00000000", 26914 => x"00000000", 26915 => x"00000000",
    26916 => x"00000000", 26917 => x"00000000", 26918 => x"00000000",
    26919 => x"00000000", 26920 => x"00000000", 26921 => x"00000000",
    26922 => x"00000000", 26923 => x"00000000", 26924 => x"00000000",
    26925 => x"00000000", 26926 => x"00000000", 26927 => x"00000000",
    26928 => x"00000000", 26929 => x"00000000", 26930 => x"00000000",
    26931 => x"00000000", 26932 => x"00000000", 26933 => x"00000000",
    26934 => x"00000000", 26935 => x"00000000", 26936 => x"00000000",
    26937 => x"00000000", 26938 => x"00000000", 26939 => x"00000000",
    26940 => x"00000000", 26941 => x"00000000", 26942 => x"00000000",
    26943 => x"00000000", 26944 => x"00000000", 26945 => x"00000000",
    26946 => x"00000000", 26947 => x"00000000", 26948 => x"00000000",
    26949 => x"00000000", 26950 => x"00000000", 26951 => x"00000000",
    26952 => x"00000000", 26953 => x"00000000", 26954 => x"00000000",
    26955 => x"00000000", 26956 => x"00000000", 26957 => x"00000000",
    26958 => x"00000000", 26959 => x"00000000", 26960 => x"00000000",
    26961 => x"00000000", 26962 => x"00000000", 26963 => x"00000000",
    26964 => x"00000000", 26965 => x"00000000", 26966 => x"00000000",
    26967 => x"00000000", 26968 => x"00000000", 26969 => x"00000000",
    26970 => x"00000000", 26971 => x"00000000", 26972 => x"00000000",
    26973 => x"00000000", 26974 => x"00000000", 26975 => x"00000000",
    26976 => x"00000000", 26977 => x"00000000", 26978 => x"00000000",
    26979 => x"00000000", 26980 => x"00000000", 26981 => x"00000000",
    26982 => x"00000000", 26983 => x"00000000", 26984 => x"00000000",
    26985 => x"00000000", 26986 => x"00000000", 26987 => x"00000000",
    26988 => x"00000000", 26989 => x"00000000", 26990 => x"00000000",
    26991 => x"00000000", 26992 => x"00000000", 26993 => x"00000000",
    26994 => x"00000000", 26995 => x"00000000", 26996 => x"00000000",
    26997 => x"00000000", 26998 => x"00000000", 26999 => x"00000000",
    27000 => x"00000000", 27001 => x"00000000", 27002 => x"00000000",
    27003 => x"00000000", 27004 => x"00000000", 27005 => x"00000000",
    27006 => x"00000000", 27007 => x"00000000", 27008 => x"00000000",
    27009 => x"00000000", 27010 => x"00000000", 27011 => x"00000000",
    27012 => x"00000000", 27013 => x"00000000", 27014 => x"00000000",
    27015 => x"00000000", 27016 => x"00000000", 27017 => x"00000000",
    27018 => x"00000000", 27019 => x"00000000", 27020 => x"00000000",
    27021 => x"00000000", 27022 => x"00000000", 27023 => x"00000000",
    27024 => x"00000000", 27025 => x"00000000", 27026 => x"00000000",
    27027 => x"00000000", 27028 => x"00000000", 27029 => x"00000000",
    27030 => x"00000000", 27031 => x"00000000", 27032 => x"00000000",
    27033 => x"00000000", 27034 => x"00000000", 27035 => x"00000000",
    27036 => x"00000000", 27037 => x"00000000", 27038 => x"00000000",
    27039 => x"00000000", 27040 => x"00000000", 27041 => x"00000000",
    27042 => x"00000000", 27043 => x"00000000", 27044 => x"00000000",
    27045 => x"00000000", 27046 => x"00000000", 27047 => x"00000000",
    27048 => x"00000000", 27049 => x"00000000", 27050 => x"00000000",
    27051 => x"00000000", 27052 => x"00000000", 27053 => x"00000000",
    27054 => x"00000000", 27055 => x"00000000", 27056 => x"00000000",
    27057 => x"00000000", 27058 => x"00000000", 27059 => x"00000000",
    27060 => x"00000000", 27061 => x"00000000", 27062 => x"00000000",
    27063 => x"00000000", 27064 => x"00000000", 27065 => x"00000000",
    27066 => x"00000000", 27067 => x"00000000", 27068 => x"00000000",
    27069 => x"00000000", 27070 => x"00000000", 27071 => x"00000000",
    27072 => x"00000000", 27073 => x"00000000", 27074 => x"00000000",
    27075 => x"00000000", 27076 => x"00000000", 27077 => x"00000000",
    27078 => x"00000000", 27079 => x"00000000", 27080 => x"00000000",
    27081 => x"00000000", 27082 => x"00000000", 27083 => x"00000000",
    27084 => x"00000000", 27085 => x"00000000", 27086 => x"00000000",
    27087 => x"00000000", 27088 => x"00000000", 27089 => x"00000000",
    27090 => x"00000000", 27091 => x"00000000", 27092 => x"00000000",
    27093 => x"00000000", 27094 => x"00000000", 27095 => x"00000000",
    27096 => x"00000000", 27097 => x"00000000", 27098 => x"00000000",
    27099 => x"00000000", 27100 => x"00000000", 27101 => x"00000000",
    27102 => x"00000000", 27103 => x"00000000", 27104 => x"00000000",
    27105 => x"00000000", 27106 => x"00000000", 27107 => x"00000000",
    27108 => x"00000000", 27109 => x"00000000", 27110 => x"00000000",
    27111 => x"00000000", 27112 => x"00000000", 27113 => x"00000000",
    27114 => x"00000000", 27115 => x"00000000", 27116 => x"00000000",
    27117 => x"00000000", 27118 => x"00000000", 27119 => x"00000000",
    27120 => x"00000000", 27121 => x"00000000", 27122 => x"00000000",
    27123 => x"00000000", 27124 => x"00000000", 27125 => x"00000000",
    27126 => x"00000000", 27127 => x"00000000", 27128 => x"00000000",
    27129 => x"00000000", 27130 => x"00000000", 27131 => x"00000000",
    27132 => x"00000000", 27133 => x"00000000", 27134 => x"00000000",
    27135 => x"00000000", 27136 => x"00000000", 27137 => x"00000000",
    27138 => x"00000000", 27139 => x"00000000", 27140 => x"00000000",
    27141 => x"00000000", 27142 => x"00000000", 27143 => x"00000000",
    27144 => x"00000000", 27145 => x"00000000", 27146 => x"00000000",
    27147 => x"00000000", 27148 => x"00000000", 27149 => x"00000000",
    27150 => x"00000000", 27151 => x"00000000", 27152 => x"00000000",
    27153 => x"00000000", 27154 => x"00000000", 27155 => x"00000000",
    27156 => x"00000000", 27157 => x"00000000", 27158 => x"00000000",
    27159 => x"00000000", 27160 => x"00000000", 27161 => x"00000000",
    27162 => x"00000000", 27163 => x"00000000", 27164 => x"00000000",
    27165 => x"00000000", 27166 => x"00000000", 27167 => x"00000000",
    27168 => x"00000000", 27169 => x"00000000", 27170 => x"00000000",
    27171 => x"00000000", 27172 => x"00000000", 27173 => x"00000000",
    27174 => x"00000000", 27175 => x"00000000", 27176 => x"00000000",
    27177 => x"00000000", 27178 => x"00000000", 27179 => x"00000000",
    27180 => x"00000000", 27181 => x"00000000", 27182 => x"00000000",
    27183 => x"00000000", 27184 => x"00000000", 27185 => x"00000000",
    27186 => x"00000000", 27187 => x"00000000", 27188 => x"00000000",
    27189 => x"00000000", 27190 => x"00000000", 27191 => x"00000000",
    27192 => x"00000000", 27193 => x"00000000", 27194 => x"00000000",
    27195 => x"00000000", 27196 => x"00000000", 27197 => x"00000000",
    27198 => x"00000000", 27199 => x"00000000", 27200 => x"00000000",
    27201 => x"00000000", 27202 => x"00000000", 27203 => x"00000000",
    27204 => x"00000000", 27205 => x"00000000", 27206 => x"00000000",
    27207 => x"00000000", 27208 => x"00000000", 27209 => x"00000000",
    27210 => x"00000000", 27211 => x"00000000", 27212 => x"00000000",
    27213 => x"00000000", 27214 => x"00000000", 27215 => x"00000000",
    27216 => x"00000000", 27217 => x"00000000", 27218 => x"00000000",
    27219 => x"00000000", 27220 => x"00000000", 27221 => x"00000000",
    27222 => x"00000000", 27223 => x"00000000", 27224 => x"00000000",
    27225 => x"00000000", 27226 => x"00000000", 27227 => x"00000000",
    27228 => x"00000000", 27229 => x"00000000", 27230 => x"00000000",
    27231 => x"00000000", 27232 => x"00000000", 27233 => x"00000000",
    27234 => x"00000000", 27235 => x"00000000", 27236 => x"00000000",
    27237 => x"00000000", 27238 => x"00000000", 27239 => x"00000000",
    27240 => x"00000000", 27241 => x"00000000", 27242 => x"00000000",
    27243 => x"00000000", 27244 => x"00000000", 27245 => x"00000000",
    27246 => x"00000000", 27247 => x"00000000", 27248 => x"00000000",
    27249 => x"00000000", 27250 => x"00000000", 27251 => x"00000000",
    27252 => x"00000000", 27253 => x"00000000", 27254 => x"00000000",
    27255 => x"00000000", 27256 => x"00000000", 27257 => x"00000000",
    27258 => x"00000000", 27259 => x"00000000", 27260 => x"00000000",
    27261 => x"00000000", 27262 => x"00000000", 27263 => x"00000000",
    27264 => x"00000000", 27265 => x"00000000", 27266 => x"00000000",
    27267 => x"00000000", 27268 => x"00000000", 27269 => x"00000000",
    27270 => x"00000000", 27271 => x"00000000", 27272 => x"00000000",
    27273 => x"00000000", 27274 => x"00000000", 27275 => x"00000000",
    27276 => x"00000000", 27277 => x"00000000", 27278 => x"00000000",
    27279 => x"00000000", 27280 => x"00000000", 27281 => x"00000000",
    27282 => x"00000000", 27283 => x"00000000", 27284 => x"00000000",
    27285 => x"00000000", 27286 => x"00000000", 27287 => x"00000000",
    27288 => x"00000000", 27289 => x"00000000", 27290 => x"00000000",
    27291 => x"00000000", 27292 => x"00000000", 27293 => x"00000000",
    27294 => x"00000000", 27295 => x"00000000", 27296 => x"00000000",
    27297 => x"00000000", 27298 => x"00000000", 27299 => x"00000000",
    27300 => x"00000000", 27301 => x"00000000", 27302 => x"00000000",
    27303 => x"00000000", 27304 => x"00000000", 27305 => x"00000000",
    27306 => x"00000000", 27307 => x"00000000", 27308 => x"00000000",
    27309 => x"00000000", 27310 => x"00000000", 27311 => x"00000000",
    27312 => x"00000000", 27313 => x"00000000", 27314 => x"00000000",
    27315 => x"00000000", 27316 => x"00000000", 27317 => x"00000000",
    27318 => x"00000000", 27319 => x"00000000", 27320 => x"00000000",
    27321 => x"00000000", 27322 => x"00000000", 27323 => x"00000000",
    27324 => x"00000000", 27325 => x"00000000", 27326 => x"00000000",
    27327 => x"00000000", 27328 => x"00000000", 27329 => x"00000000",
    27330 => x"00000000", 27331 => x"00000000", 27332 => x"00000000",
    27333 => x"00000000", 27334 => x"00000000", 27335 => x"00000000",
    27336 => x"00000000", 27337 => x"00000000", 27338 => x"00000000",
    27339 => x"00000000", 27340 => x"00000000", 27341 => x"00000000",
    27342 => x"00000000", 27343 => x"00000000", 27344 => x"00000000",
    27345 => x"00000000", 27346 => x"00000000", 27347 => x"00000000",
    27348 => x"00000000", 27349 => x"00000000", 27350 => x"00000000",
    27351 => x"00000000", 27352 => x"00000000", 27353 => x"00000000",
    27354 => x"00000000", 27355 => x"00000000", 27356 => x"00000000",
    27357 => x"00000000", 27358 => x"00000000", 27359 => x"00000000",
    27360 => x"00000000", 27361 => x"00000000", 27362 => x"00000000",
    27363 => x"00000000", 27364 => x"00000000", 27365 => x"00000000",
    27366 => x"00000000", 27367 => x"00000000", 27368 => x"00000000",
    27369 => x"00000000", 27370 => x"00000000", 27371 => x"00000000",
    27372 => x"00000000", 27373 => x"00000000", 27374 => x"00000000",
    27375 => x"00000000", 27376 => x"00000000", 27377 => x"00000000",
    27378 => x"00000000", 27379 => x"00000000", 27380 => x"00000000",
    27381 => x"00000000", 27382 => x"00000000", 27383 => x"00000000",
    27384 => x"00000000", 27385 => x"00000000", 27386 => x"00000000",
    27387 => x"00000000", 27388 => x"00000000", 27389 => x"00000000",
    27390 => x"00000000", 27391 => x"00000000", 27392 => x"00000000",
    27393 => x"00000000", 27394 => x"00000000", 27395 => x"00000000",
    27396 => x"00000000", 27397 => x"00000000", 27398 => x"00000000",
    27399 => x"00000000", 27400 => x"00000000", 27401 => x"00000000",
    27402 => x"00000000", 27403 => x"00000000", 27404 => x"00000000",
    27405 => x"00000000", 27406 => x"00000000", 27407 => x"00000000",
    27408 => x"00000000", 27409 => x"00000000", 27410 => x"00000000",
    27411 => x"00000000", 27412 => x"00000000", 27413 => x"00000000",
    27414 => x"00000000", 27415 => x"00000000", 27416 => x"00000000",
    27417 => x"00000000", 27418 => x"00000000", 27419 => x"00000000",
    27420 => x"00000000", 27421 => x"00000000", 27422 => x"00000000",
    27423 => x"00000000", 27424 => x"00000000", 27425 => x"00000000",
    27426 => x"00000000", 27427 => x"00000000", 27428 => x"00000000",
    27429 => x"00000000", 27430 => x"00000000", 27431 => x"00000000",
    27432 => x"00000000", 27433 => x"00000000", 27434 => x"00000000",
    27435 => x"00000000", 27436 => x"00000000", 27437 => x"00000000",
    27438 => x"00000000", 27439 => x"00000000", 27440 => x"00000000",
    27441 => x"00000000", 27442 => x"00000000", 27443 => x"00000000",
    27444 => x"00000000", 27445 => x"00000000", 27446 => x"00000000",
    27447 => x"00000000", 27448 => x"00000000", 27449 => x"00000000",
    27450 => x"00000000", 27451 => x"00000000", 27452 => x"00000000",
    27453 => x"00000000", 27454 => x"00000000", 27455 => x"00000000",
    27456 => x"00000000", 27457 => x"00000000", 27458 => x"00000000",
    27459 => x"00000000", 27460 => x"00000000", 27461 => x"00000000",
    27462 => x"00000000", 27463 => x"00000000", 27464 => x"00000000",
    27465 => x"00000000", 27466 => x"00000000", 27467 => x"00000000",
    27468 => x"00000000", 27469 => x"00000000", 27470 => x"00000000",
    27471 => x"00000000", 27472 => x"00000000", 27473 => x"00000000",
    27474 => x"00000000", 27475 => x"00000000", 27476 => x"00000000",
    27477 => x"00000000", 27478 => x"00000000", 27479 => x"00000000",
    27480 => x"00000000", 27481 => x"00000000", 27482 => x"00000000",
    27483 => x"00000000", 27484 => x"00000000", 27485 => x"00000000",
    27486 => x"00000000", 27487 => x"00000000", 27488 => x"00000000",
    27489 => x"00000000", 27490 => x"00000000", 27491 => x"00000000",
    27492 => x"00000000", 27493 => x"00000000", 27494 => x"00000000",
    27495 => x"00000000", 27496 => x"00000000", 27497 => x"00000000",
    27498 => x"00000000", 27499 => x"00000000", 27500 => x"00000000",
    27501 => x"00000000", 27502 => x"00000000", 27503 => x"00000000",
    27504 => x"00000000", 27505 => x"00000000", 27506 => x"00000000",
    27507 => x"00000000", 27508 => x"00000000", 27509 => x"00000000",
    27510 => x"00000000", 27511 => x"00000000", 27512 => x"00000000",
    27513 => x"00000000", 27514 => x"00000000", 27515 => x"00000000",
    27516 => x"00000000", 27517 => x"00000000", 27518 => x"00000000",
    27519 => x"00000000", 27520 => x"00000000", 27521 => x"00000000",
    27522 => x"00000000", 27523 => x"00000000", 27524 => x"00000000",
    27525 => x"00000000", 27526 => x"00000000", 27527 => x"00000000",
    27528 => x"00000000", 27529 => x"00000000", 27530 => x"00000000",
    27531 => x"00000000", 27532 => x"00000000", 27533 => x"00000000",
    27534 => x"00000000", 27535 => x"00000000", 27536 => x"00000000",
    27537 => x"00000000", 27538 => x"00000000", 27539 => x"00000000",
    27540 => x"00000000", 27541 => x"00000000", 27542 => x"00000000",
    27543 => x"00000000", 27544 => x"00000000", 27545 => x"00000000",
    27546 => x"00000000", 27547 => x"00000000", 27548 => x"00000000",
    27549 => x"00000000", 27550 => x"00000000", 27551 => x"00000000",
    27552 => x"00000000", 27553 => x"00000000", 27554 => x"00000000",
    27555 => x"00000000", 27556 => x"00000000", 27557 => x"00000000",
    27558 => x"00000000", 27559 => x"00000000", 27560 => x"00000000",
    27561 => x"00000000", 27562 => x"00000000", 27563 => x"00000000",
    27564 => x"00000000", 27565 => x"00000000", 27566 => x"00000000",
    27567 => x"00000000", 27568 => x"00000000", 27569 => x"00000000",
    27570 => x"00000000", 27571 => x"00000000", 27572 => x"00000000",
    27573 => x"00000000", 27574 => x"00000000", 27575 => x"00000000",
    27576 => x"00000000", 27577 => x"00000000", 27578 => x"00000000",
    27579 => x"00000000", 27580 => x"00000000", 27581 => x"00000000",
    27582 => x"00000000", 27583 => x"00000000", 27584 => x"00000000",
    27585 => x"00000000", 27586 => x"00000000", 27587 => x"00000000",
    27588 => x"00000000", 27589 => x"00000000", 27590 => x"00000000",
    27591 => x"00000000", 27592 => x"00000000", 27593 => x"00000000",
    27594 => x"00000000", 27595 => x"00000000", 27596 => x"00000000",
    27597 => x"00000000", 27598 => x"00000000", 27599 => x"00000000",
    27600 => x"00000000", 27601 => x"00000000", 27602 => x"00000000",
    27603 => x"00000000", 27604 => x"00000000", 27605 => x"00000000",
    27606 => x"00000000", 27607 => x"00000000", 27608 => x"00000000",
    27609 => x"00000000", 27610 => x"00000000", 27611 => x"00000000",
    27612 => x"00000000", 27613 => x"00000000", 27614 => x"00000000",
    27615 => x"00000000", 27616 => x"00000000", 27617 => x"00000000",
    27618 => x"00000000", 27619 => x"00000000", 27620 => x"00000000",
    27621 => x"00000000", 27622 => x"00000000", 27623 => x"00000000",
    27624 => x"00000000", 27625 => x"00000000", 27626 => x"00000000",
    27627 => x"00000000", 27628 => x"00000000", 27629 => x"00000000",
    27630 => x"00000000", 27631 => x"00000000", 27632 => x"00000000",
    27633 => x"00000000", 27634 => x"00000000", 27635 => x"00000000",
    27636 => x"00000000", 27637 => x"00000000", 27638 => x"00000000",
    27639 => x"00000000", 27640 => x"00000000", 27641 => x"00000000",
    27642 => x"00000000", 27643 => x"00000000", 27644 => x"00000000",
    27645 => x"00000000", 27646 => x"00000000", 27647 => x"00000000",
    27648 => x"00000000", 27649 => x"00000000", 27650 => x"00000000",
    27651 => x"00000000", 27652 => x"00000000", 27653 => x"00000000",
    27654 => x"00000000", 27655 => x"00000000", 27656 => x"00000000",
    27657 => x"00000000", 27658 => x"00000000", 27659 => x"00000000",
    27660 => x"00000000", 27661 => x"00000000", 27662 => x"00000000",
    27663 => x"00000000", 27664 => x"00000000", 27665 => x"00000000",
    27666 => x"00000000", 27667 => x"00000000", 27668 => x"00000000",
    27669 => x"00000000", 27670 => x"00000000", 27671 => x"00000000",
    27672 => x"00000000", 27673 => x"00000000", 27674 => x"00000000",
    27675 => x"00000000", 27676 => x"00000000", 27677 => x"00000000",
    27678 => x"00000000", 27679 => x"00000000", 27680 => x"00000000",
    27681 => x"00000000", 27682 => x"00000000", 27683 => x"00000000",
    27684 => x"00000000", 27685 => x"00000000", 27686 => x"00000000",
    27687 => x"00000000", 27688 => x"00000000", 27689 => x"00000000",
    27690 => x"00000000", 27691 => x"00000000", 27692 => x"00000000",
    27693 => x"00000000", 27694 => x"00000000", 27695 => x"00000000",
    27696 => x"00000000", 27697 => x"00000000", 27698 => x"00000000",
    27699 => x"00000000", 27700 => x"00000000", 27701 => x"00000000",
    27702 => x"00000000", 27703 => x"00000000", 27704 => x"00000000",
    27705 => x"00000000", 27706 => x"00000000", 27707 => x"00000000",
    27708 => x"00000000", 27709 => x"00000000", 27710 => x"00000000",
    27711 => x"00000000", 27712 => x"00000000", 27713 => x"00000000",
    27714 => x"00000000", 27715 => x"00000000", 27716 => x"00000000",
    27717 => x"00000000", 27718 => x"00000000", 27719 => x"00000000",
    27720 => x"00000000", 27721 => x"00000000", 27722 => x"00000000",
    27723 => x"00000000", 27724 => x"00000000", 27725 => x"00000000",
    27726 => x"00000000", 27727 => x"00000000", 27728 => x"00000000",
    27729 => x"00000000", 27730 => x"00000000", 27731 => x"00000000",
    27732 => x"00000000", 27733 => x"00000000", 27734 => x"00000000",
    27735 => x"00000000", 27736 => x"00000000", 27737 => x"00000000",
    27738 => x"00000000", 27739 => x"00000000", 27740 => x"00000000",
    27741 => x"00000000", 27742 => x"00000000", 27743 => x"00000000",
    27744 => x"00000000", 27745 => x"00000000", 27746 => x"00000000",
    27747 => x"00000000", 27748 => x"00000000", 27749 => x"00000000",
    27750 => x"00000000", 27751 => x"00000000", 27752 => x"00000000",
    27753 => x"00000000", 27754 => x"00000000", 27755 => x"00000000",
    27756 => x"00000000", 27757 => x"00000000", 27758 => x"00000000",
    27759 => x"00000000", 27760 => x"00000000", 27761 => x"00000000",
    27762 => x"00000000", 27763 => x"00000000", 27764 => x"00000000",
    27765 => x"00000000", 27766 => x"00000000", 27767 => x"00000000",
    27768 => x"00000000", 27769 => x"00000000", 27770 => x"00000000",
    27771 => x"00000000", 27772 => x"00000000", 27773 => x"00000000",
    27774 => x"00000000", 27775 => x"00000000", 27776 => x"00000000",
    27777 => x"00000000", 27778 => x"00000000", 27779 => x"00000000",
    27780 => x"00000000", 27781 => x"00000000", 27782 => x"00000000",
    27783 => x"00000000", 27784 => x"00000000", 27785 => x"00000000",
    27786 => x"00000000", 27787 => x"00000000", 27788 => x"00000000",
    27789 => x"00000000", 27790 => x"00000000", 27791 => x"00000000",
    27792 => x"00000000", 27793 => x"00000000", 27794 => x"00000000",
    27795 => x"00000000", 27796 => x"00000000", 27797 => x"00000000",
    27798 => x"00000000", 27799 => x"00000000", 27800 => x"00000000",
    27801 => x"00000000", 27802 => x"00000000", 27803 => x"00000000",
    27804 => x"00000000", 27805 => x"00000000", 27806 => x"00000000",
    27807 => x"00000000", 27808 => x"00000000", 27809 => x"00000000",
    27810 => x"00000000", 27811 => x"00000000", 27812 => x"00000000",
    27813 => x"00000000", 27814 => x"00000000", 27815 => x"00000000",
    27816 => x"00000000", 27817 => x"00000000", 27818 => x"00000000",
    27819 => x"00000000", 27820 => x"00000000", 27821 => x"00000000",
    27822 => x"00000000", 27823 => x"00000000", 27824 => x"00000000",
    27825 => x"00000000", 27826 => x"00000000", 27827 => x"00000000",
    27828 => x"00000000", 27829 => x"00000000", 27830 => x"00000000",
    27831 => x"00000000", 27832 => x"00000000", 27833 => x"00000000",
    27834 => x"00000000", 27835 => x"00000000", 27836 => x"00000000",
    27837 => x"00000000", 27838 => x"00000000", 27839 => x"00000000",
    27840 => x"00000000", 27841 => x"00000000", 27842 => x"00000000",
    27843 => x"00000000", 27844 => x"00000000", 27845 => x"00000000",
    27846 => x"00000000", 27847 => x"00000000", 27848 => x"00000000",
    27849 => x"00000000", 27850 => x"00000000", 27851 => x"00000000",
    27852 => x"00000000", 27853 => x"00000000", 27854 => x"00000000",
    27855 => x"00000000", 27856 => x"00000000", 27857 => x"00000000",
    27858 => x"00000000", 27859 => x"00000000", 27860 => x"00000000",
    27861 => x"00000000", 27862 => x"00000000", 27863 => x"00000000",
    27864 => x"00000000", 27865 => x"00000000", 27866 => x"00000000",
    27867 => x"00000000", 27868 => x"00000000", 27869 => x"00000000",
    27870 => x"00000000", 27871 => x"00000000", 27872 => x"00000000",
    27873 => x"00000000", 27874 => x"00000000", 27875 => x"00000000",
    27876 => x"00000000", 27877 => x"00000000", 27878 => x"00000000",
    27879 => x"00000000", 27880 => x"00000000", 27881 => x"00000000",
    27882 => x"00000000", 27883 => x"00000000", 27884 => x"00000000",
    27885 => x"00000000", 27886 => x"00000000", 27887 => x"00000000",
    27888 => x"00000000", 27889 => x"00000000", 27890 => x"00000000",
    27891 => x"00000000", 27892 => x"00000000", 27893 => x"00000000",
    27894 => x"00000000", 27895 => x"00000000", 27896 => x"00000000",
    27897 => x"00000000", 27898 => x"00000000", 27899 => x"00000000",
    27900 => x"00000000", 27901 => x"00000000", 27902 => x"00000000",
    27903 => x"00000000", 27904 => x"00000000", 27905 => x"00000000",
    27906 => x"00000000", 27907 => x"00000000", 27908 => x"00000000",
    27909 => x"00000000", 27910 => x"00000000", 27911 => x"00000000",
    27912 => x"00000000", 27913 => x"00000000", 27914 => x"00000000",
    27915 => x"00000000", 27916 => x"00000000", 27917 => x"00000000",
    27918 => x"00000000", 27919 => x"00000000", 27920 => x"00000000",
    27921 => x"00000000", 27922 => x"00000000", 27923 => x"00000000",
    27924 => x"00000000", 27925 => x"00000000", 27926 => x"00000000",
    27927 => x"00000000", 27928 => x"00000000", 27929 => x"00000000",
    27930 => x"00000000", 27931 => x"00000000", 27932 => x"00000000",
    27933 => x"00000000", 27934 => x"00000000", 27935 => x"00000000",
    27936 => x"00000000", 27937 => x"00000000", 27938 => x"00000000",
    27939 => x"00000000", 27940 => x"00000000", 27941 => x"00000000",
    27942 => x"00000000", 27943 => x"00000000", 27944 => x"00000000",
    27945 => x"00000000", 27946 => x"00000000", 27947 => x"00000000",
    27948 => x"00000000", 27949 => x"00000000", 27950 => x"00000000",
    27951 => x"00000000", 27952 => x"00000000", 27953 => x"00000000",
    27954 => x"00000000", 27955 => x"00000000", 27956 => x"00000000",
    27957 => x"00000000", 27958 => x"00000000", 27959 => x"00000000",
    27960 => x"00000000", 27961 => x"00000000", 27962 => x"00000000",
    27963 => x"00000000", 27964 => x"00000000", 27965 => x"00000000",
    27966 => x"00000000", 27967 => x"00000000", 27968 => x"00000000",
    27969 => x"00000000", 27970 => x"00000000", 27971 => x"00000000",
    27972 => x"00000000", 27973 => x"00000000", 27974 => x"00000000",
    27975 => x"00000000", 27976 => x"00000000", 27977 => x"00000000",
    27978 => x"00000000", 27979 => x"00000000", 27980 => x"00000000",
    27981 => x"00000000", 27982 => x"00000000", 27983 => x"00000000",
    27984 => x"00000000", 27985 => x"00000000", 27986 => x"00000000",
    27987 => x"00000000", 27988 => x"00000000", 27989 => x"00000000",
    27990 => x"00000000", 27991 => x"00000000", 27992 => x"00000000",
    27993 => x"00000000", 27994 => x"00000000", 27995 => x"00000000",
    27996 => x"00000000", 27997 => x"00000000", 27998 => x"00000000",
    27999 => x"00000000", 28000 => x"00000000", 28001 => x"00000000",
    28002 => x"00000000", 28003 => x"00000000", 28004 => x"00000000",
    28005 => x"00000000", 28006 => x"00000000", 28007 => x"00000000",
    28008 => x"00000000", 28009 => x"00000000", 28010 => x"00000000",
    28011 => x"00000000", 28012 => x"00000000", 28013 => x"00000000",
    28014 => x"00000000", 28015 => x"00000000", 28016 => x"00000000",
    28017 => x"00000000", 28018 => x"00000000", 28019 => x"00000000",
    28020 => x"00000000", 28021 => x"00000000", 28022 => x"00000000",
    28023 => x"00000000", 28024 => x"00000000", 28025 => x"00000000",
    28026 => x"00000000", 28027 => x"00000000", 28028 => x"00000000",
    28029 => x"00000000", 28030 => x"00000000", 28031 => x"00000000",
    28032 => x"00000000", 28033 => x"00000000", 28034 => x"00000000",
    28035 => x"00000000", 28036 => x"00000000", 28037 => x"00000000",
    28038 => x"00000000", 28039 => x"00000000", 28040 => x"00000000",
    28041 => x"00000000", 28042 => x"00000000", 28043 => x"00000000",
    28044 => x"00000000", 28045 => x"00000000", 28046 => x"00000000",
    28047 => x"00000000", 28048 => x"00000000", 28049 => x"00000000",
    28050 => x"00000000", 28051 => x"00000000", 28052 => x"00000000",
    28053 => x"00000000", 28054 => x"00000000", 28055 => x"00000000",
    28056 => x"00000000", 28057 => x"00000000", 28058 => x"00000000",
    28059 => x"00000000", 28060 => x"00000000", 28061 => x"00000000",
    28062 => x"00000000", 28063 => x"00000000", 28064 => x"00000000",
    28065 => x"00000000", 28066 => x"00000000", 28067 => x"00000000",
    28068 => x"00000000", 28069 => x"00000000", 28070 => x"00000000",
    28071 => x"00000000", 28072 => x"00000000", 28073 => x"00000000",
    28074 => x"00000000", 28075 => x"00000000", 28076 => x"00000000",
    28077 => x"00000000", 28078 => x"00000000", 28079 => x"00000000",
    28080 => x"00000000", 28081 => x"00000000", 28082 => x"00000000",
    28083 => x"00000000", 28084 => x"00000000", 28085 => x"00000000",
    28086 => x"00000000", 28087 => x"00000000", 28088 => x"00000000",
    28089 => x"00000000", 28090 => x"00000000", 28091 => x"00000000",
    28092 => x"00000000", 28093 => x"00000000", 28094 => x"00000000",
    28095 => x"00000000", 28096 => x"00000000", 28097 => x"00000000",
    28098 => x"00000000", 28099 => x"00000000", 28100 => x"00000000",
    28101 => x"00000000", 28102 => x"00000000", 28103 => x"00000000",
    28104 => x"00000000", 28105 => x"00000000", 28106 => x"00000000",
    28107 => x"00000000", 28108 => x"00000000", 28109 => x"00000000",
    28110 => x"00000000", 28111 => x"00000000", 28112 => x"00000000",
    28113 => x"00000000", 28114 => x"00000000", 28115 => x"00000000",
    28116 => x"00000000", 28117 => x"00000000", 28118 => x"00000000",
    28119 => x"00000000", 28120 => x"00000000", 28121 => x"00000000",
    28122 => x"00000000", 28123 => x"00000000", 28124 => x"00000000",
    28125 => x"00000000", 28126 => x"00000000", 28127 => x"00000000",
    28128 => x"00000000", 28129 => x"00000000", 28130 => x"00000000",
    28131 => x"00000000", 28132 => x"00000000", 28133 => x"00000000",
    28134 => x"00000000", 28135 => x"00000000", 28136 => x"00000000",
    28137 => x"00000000", 28138 => x"00000000", 28139 => x"00000000",
    28140 => x"00000000", 28141 => x"00000000", 28142 => x"00000000",
    28143 => x"00000000", 28144 => x"00000000", 28145 => x"00000000",
    28146 => x"00000000", 28147 => x"00000000", 28148 => x"00000000",
    28149 => x"00000000", 28150 => x"00000000", 28151 => x"00000000",
    28152 => x"00000000", 28153 => x"00000000", 28154 => x"00000000",
    28155 => x"00000000", 28156 => x"00000000", 28157 => x"00000000",
    28158 => x"00000000", 28159 => x"00000000", 28160 => x"00000000",
    28161 => x"00000000", 28162 => x"00000000", 28163 => x"00000000",
    28164 => x"00000000", 28165 => x"00000000", 28166 => x"00000000",
    28167 => x"00000000", 28168 => x"00000000", 28169 => x"00000000",
    28170 => x"00000000", 28171 => x"00000000", 28172 => x"00000000",
    28173 => x"00000000", 28174 => x"00000000", 28175 => x"00000000",
    28176 => x"00000000", 28177 => x"00000000", 28178 => x"00000000",
    28179 => x"00000000", 28180 => x"00000000", 28181 => x"00000000",
    28182 => x"00000000", 28183 => x"00000000", 28184 => x"00000000",
    28185 => x"00000000", 28186 => x"00000000", 28187 => x"00000000",
    28188 => x"00000000", 28189 => x"00000000", 28190 => x"00000000",
    28191 => x"00000000", 28192 => x"00000000", 28193 => x"00000000",
    28194 => x"00000000", 28195 => x"00000000", 28196 => x"00000000",
    28197 => x"00000000", 28198 => x"00000000", 28199 => x"00000000",
    28200 => x"00000000", 28201 => x"00000000", 28202 => x"00000000",
    28203 => x"00000000", 28204 => x"00000000", 28205 => x"00000000",
    28206 => x"00000000", 28207 => x"00000000", 28208 => x"00000000",
    28209 => x"00000000", 28210 => x"00000000", 28211 => x"00000000",
    28212 => x"00000000", 28213 => x"00000000", 28214 => x"00000000",
    28215 => x"00000000", 28216 => x"00000000", 28217 => x"00000000",
    28218 => x"00000000", 28219 => x"00000000", 28220 => x"00000000",
    28221 => x"00000000", 28222 => x"00000000", 28223 => x"00000000",
    28224 => x"00000000", 28225 => x"00000000", 28226 => x"00000000",
    28227 => x"00000000", 28228 => x"00000000", 28229 => x"00000000",
    28230 => x"00000000", 28231 => x"00000000", 28232 => x"00000000",
    28233 => x"00000000", 28234 => x"00000000", 28235 => x"00000000",
    28236 => x"00000000", 28237 => x"00000000", 28238 => x"00000000",
    28239 => x"00000000", 28240 => x"00000000", 28241 => x"00000000",
    28242 => x"00000000", 28243 => x"00000000", 28244 => x"00000000",
    28245 => x"00000000", 28246 => x"00000000", 28247 => x"00000000",
    28248 => x"00000000", 28249 => x"00000000", 28250 => x"00000000",
    28251 => x"00000000", 28252 => x"00000000", 28253 => x"00000000",
    28254 => x"00000000", 28255 => x"00000000", 28256 => x"00000000",
    28257 => x"00000000", 28258 => x"00000000", 28259 => x"00000000",
    28260 => x"00000000", 28261 => x"00000000", 28262 => x"00000000",
    28263 => x"00000000", 28264 => x"00000000", 28265 => x"00000000",
    28266 => x"00000000", 28267 => x"00000000", 28268 => x"00000000",
    28269 => x"00000000", 28270 => x"00000000", 28271 => x"00000000",
    28272 => x"00000000", 28273 => x"00000000", 28274 => x"00000000",
    28275 => x"00000000", 28276 => x"00000000", 28277 => x"00000000",
    28278 => x"00000000", 28279 => x"00000000", 28280 => x"00000000",
    28281 => x"00000000", 28282 => x"00000000", 28283 => x"00000000",
    28284 => x"00000000", 28285 => x"00000000", 28286 => x"00000000",
    28287 => x"00000000", 28288 => x"00000000", 28289 => x"00000000",
    28290 => x"00000000", 28291 => x"00000000", 28292 => x"00000000",
    28293 => x"00000000", 28294 => x"00000000", 28295 => x"00000000",
    28296 => x"00000000", 28297 => x"00000000", 28298 => x"00000000",
    28299 => x"00000000", 28300 => x"00000000", 28301 => x"00000000",
    28302 => x"00000000", 28303 => x"00000000", 28304 => x"00000000",
    28305 => x"00000000", 28306 => x"00000000", 28307 => x"00000000",
    28308 => x"00000000", 28309 => x"00000000", 28310 => x"00000000",
    28311 => x"00000000", 28312 => x"00000000", 28313 => x"00000000",
    28314 => x"00000000", 28315 => x"00000000", 28316 => x"00000000",
    28317 => x"00000000", 28318 => x"00000000", 28319 => x"00000000",
    28320 => x"00000000", 28321 => x"00000000", 28322 => x"00000000",
    28323 => x"00000000", 28324 => x"00000000", 28325 => x"00000000",
    28326 => x"00000000", 28327 => x"00000000", 28328 => x"00000000",
    28329 => x"00000000", 28330 => x"00000000", 28331 => x"00000000",
    28332 => x"00000000", 28333 => x"00000000", 28334 => x"00000000",
    28335 => x"00000000", 28336 => x"00000000", 28337 => x"00000000",
    28338 => x"00000000", 28339 => x"00000000", 28340 => x"00000000",
    28341 => x"00000000", 28342 => x"00000000", 28343 => x"00000000",
    28344 => x"00000000", 28345 => x"00000000", 28346 => x"00000000",
    28347 => x"00000000", 28348 => x"00000000", 28349 => x"00000000",
    28350 => x"00000000", 28351 => x"00000000", 28352 => x"00000000",
    28353 => x"00000000", 28354 => x"00000000", 28355 => x"00000000",
    28356 => x"00000000", 28357 => x"00000000", 28358 => x"00000000",
    28359 => x"00000000", 28360 => x"00000000", 28361 => x"00000000",
    28362 => x"00000000", 28363 => x"00000000", 28364 => x"00000000",
    28365 => x"00000000", 28366 => x"00000000", 28367 => x"00000000",
    28368 => x"00000000", 28369 => x"00000000", 28370 => x"00000000",
    28371 => x"00000000", 28372 => x"00000000", 28373 => x"00000000",
    28374 => x"00000000", 28375 => x"00000000", 28376 => x"00000000",
    28377 => x"00000000", 28378 => x"00000000", 28379 => x"00000000",
    28380 => x"00000000", 28381 => x"00000000", 28382 => x"00000000",
    28383 => x"00000000", 28384 => x"00000000", 28385 => x"00000000",
    28386 => x"00000000", 28387 => x"00000000", 28388 => x"00000000",
    28389 => x"00000000", 28390 => x"00000000", 28391 => x"00000000",
    28392 => x"00000000", 28393 => x"00000000", 28394 => x"00000000",
    28395 => x"00000000", 28396 => x"00000000", 28397 => x"00000000",
    28398 => x"00000000", 28399 => x"00000000", 28400 => x"00000000",
    28401 => x"00000000", 28402 => x"00000000", 28403 => x"00000000",
    28404 => x"00000000", 28405 => x"00000000", 28406 => x"00000000",
    28407 => x"00000000", 28408 => x"00000000", 28409 => x"00000000",
    28410 => x"00000000", 28411 => x"00000000", 28412 => x"00000000",
    28413 => x"00000000", 28414 => x"00000000", 28415 => x"00000000",
    28416 => x"00000000", 28417 => x"00000000", 28418 => x"00000000",
    28419 => x"00000000", 28420 => x"00000000", 28421 => x"00000000",
    28422 => x"00000000", 28423 => x"00000000", 28424 => x"00000000",
    28425 => x"00000000", 28426 => x"00000000", 28427 => x"00000000",
    28428 => x"00000000", 28429 => x"00000000", 28430 => x"00000000",
    28431 => x"00000000", 28432 => x"00000000", 28433 => x"00000000",
    28434 => x"00000000", 28435 => x"00000000", 28436 => x"00000000",
    28437 => x"00000000", 28438 => x"00000000", 28439 => x"00000000",
    28440 => x"00000000", 28441 => x"00000000", 28442 => x"00000000",
    28443 => x"00000000", 28444 => x"00000000", 28445 => x"00000000",
    28446 => x"00000000", 28447 => x"00000000", 28448 => x"00000000",
    28449 => x"00000000", 28450 => x"00000000", 28451 => x"00000000",
    28452 => x"00000000", 28453 => x"00000000", 28454 => x"00000000",
    28455 => x"00000000", 28456 => x"00000000", 28457 => x"00000000",
    28458 => x"00000000", 28459 => x"00000000", 28460 => x"00000000",
    28461 => x"00000000", 28462 => x"00000000", 28463 => x"00000000",
    28464 => x"00000000", 28465 => x"00000000", 28466 => x"00000000",
    28467 => x"00000000", 28468 => x"00000000", 28469 => x"00000000",
    28470 => x"00000000", 28471 => x"00000000", 28472 => x"00000000",
    28473 => x"00000000", 28474 => x"00000000", 28475 => x"00000000",
    28476 => x"00000000", 28477 => x"00000000", 28478 => x"00000000",
    28479 => x"00000000", 28480 => x"00000000", 28481 => x"00000000",
    28482 => x"00000000", 28483 => x"00000000", 28484 => x"00000000",
    28485 => x"00000000", 28486 => x"00000000", 28487 => x"00000000",
    28488 => x"00000000", 28489 => x"00000000", 28490 => x"00000000",
    28491 => x"00000000", 28492 => x"00000000", 28493 => x"00000000",
    28494 => x"00000000", 28495 => x"00000000", 28496 => x"00000000",
    28497 => x"00000000", 28498 => x"00000000", 28499 => x"00000000",
    28500 => x"00000000", 28501 => x"00000000", 28502 => x"00000000",
    28503 => x"00000000", 28504 => x"00000000", 28505 => x"00000000",
    28506 => x"00000000", 28507 => x"00000000", 28508 => x"00000000",
    28509 => x"00000000", 28510 => x"00000000", 28511 => x"00000000",
    28512 => x"00000000", 28513 => x"00000000", 28514 => x"00000000",
    28515 => x"00000000", 28516 => x"00000000", 28517 => x"00000000",
    28518 => x"00000000", 28519 => x"00000000", 28520 => x"00000000",
    28521 => x"00000000", 28522 => x"00000000", 28523 => x"00000000",
    28524 => x"00000000", 28525 => x"00000000", 28526 => x"00000000",
    28527 => x"00000000", 28528 => x"00000000", 28529 => x"00000000",
    28530 => x"00000000", 28531 => x"00000000", 28532 => x"00000000",
    28533 => x"00000000", 28534 => x"00000000", 28535 => x"00000000",
    28536 => x"00000000", 28537 => x"00000000", 28538 => x"00000000",
    28539 => x"00000000", 28540 => x"00000000", 28541 => x"00000000",
    28542 => x"00000000", 28543 => x"00000000", 28544 => x"00000000",
    28545 => x"00000000", 28546 => x"00000000", 28547 => x"00000000",
    28548 => x"00000000", 28549 => x"00000000", 28550 => x"00000000",
    28551 => x"00000000", 28552 => x"00000000", 28553 => x"00000000",
    28554 => x"00000000", 28555 => x"00000000", 28556 => x"00000000",
    28557 => x"00000000", 28558 => x"00000000", 28559 => x"00000000",
    28560 => x"00000000", 28561 => x"00000000", 28562 => x"00000000",
    28563 => x"00000000", 28564 => x"00000000", 28565 => x"00000000",
    28566 => x"00000000", 28567 => x"00000000", 28568 => x"00000000",
    28569 => x"00000000", 28570 => x"00000000", 28571 => x"00000000",
    28572 => x"00000000", 28573 => x"00000000", 28574 => x"00000000",
    28575 => x"00000000", 28576 => x"00000000", 28577 => x"00000000",
    28578 => x"00000000", 28579 => x"00000000", 28580 => x"00000000",
    28581 => x"00000000", 28582 => x"00000000", 28583 => x"00000000",
    28584 => x"00000000", 28585 => x"00000000", 28586 => x"00000000",
    28587 => x"00000000", 28588 => x"00000000", 28589 => x"00000000",
    28590 => x"00000000", 28591 => x"00000000", 28592 => x"00000000",
    28593 => x"00000000", 28594 => x"00000000", 28595 => x"00000000",
    28596 => x"00000000", 28597 => x"00000000", 28598 => x"00000000",
    28599 => x"00000000", 28600 => x"00000000", 28601 => x"00000000",
    28602 => x"00000000", 28603 => x"00000000", 28604 => x"00000000",
    28605 => x"00000000", 28606 => x"00000000", 28607 => x"00000000",
    28608 => x"00000000", 28609 => x"00000000", 28610 => x"00000000",
    28611 => x"00000000", 28612 => x"00000000", 28613 => x"00000000",
    28614 => x"00000000", 28615 => x"00000000", 28616 => x"00000000",
    28617 => x"00000000", 28618 => x"00000000", 28619 => x"00000000",
    28620 => x"00000000", 28621 => x"00000000", 28622 => x"00000000",
    28623 => x"00000000", 28624 => x"00000000", 28625 => x"00000000",
    28626 => x"00000000", 28627 => x"00000000", 28628 => x"00000000",
    28629 => x"00000000", 28630 => x"00000000", 28631 => x"00000000",
    28632 => x"00000000", 28633 => x"00000000", 28634 => x"00000000",
    28635 => x"00000000", 28636 => x"00000000", 28637 => x"00000000",
    28638 => x"00000000", 28639 => x"00000000", 28640 => x"00000000",
    28641 => x"00000000", 28642 => x"00000000", 28643 => x"00000000",
    28644 => x"00000000", 28645 => x"00000000", 28646 => x"00000000",
    28647 => x"00000000", 28648 => x"00000000", 28649 => x"00000000",
    28650 => x"00000000", 28651 => x"00000000", 28652 => x"00000000",
    28653 => x"00000000", 28654 => x"00000000", 28655 => x"00000000",
    28656 => x"00000000", 28657 => x"00000000", 28658 => x"00000000",
    28659 => x"00000000", 28660 => x"00000000", 28661 => x"00000000",
    28662 => x"00000000", 28663 => x"00000000", 28664 => x"00000000",
    28665 => x"00000000", 28666 => x"00000000", 28667 => x"00000000",
    28668 => x"00000000", 28669 => x"00000000", 28670 => x"00000000",
    28671 => x"00000000", 28672 => x"00000000", 28673 => x"00000000",
    28674 => x"00000000", 28675 => x"00000000", 28676 => x"00000000",
    28677 => x"00000000", 28678 => x"00000000", 28679 => x"00000000",
    28680 => x"00000000", 28681 => x"00000000", 28682 => x"00000000",
    28683 => x"00000000", 28684 => x"00000000", 28685 => x"00000000",
    28686 => x"00000000", 28687 => x"00000000", 28688 => x"00000000",
    28689 => x"00000000", 28690 => x"00000000", 28691 => x"00000000",
    28692 => x"00000000", 28693 => x"00000000", 28694 => x"00000000",
    28695 => x"00000000", 28696 => x"00000000", 28697 => x"00000000",
    28698 => x"00000000", 28699 => x"00000000", 28700 => x"00000000",
    28701 => x"00000000", 28702 => x"00000000", 28703 => x"00000000",
    28704 => x"00000000", 28705 => x"00000000", 28706 => x"00000000",
    28707 => x"00000000", 28708 => x"00000000", 28709 => x"00000000",
    28710 => x"00000000", 28711 => x"00000000", 28712 => x"00000000",
    28713 => x"00000000", 28714 => x"00000000", 28715 => x"00000000",
    28716 => x"00000000", 28717 => x"00000000", 28718 => x"00000000",
    28719 => x"00000000", 28720 => x"00000000", 28721 => x"00000000",
    28722 => x"00000000", 28723 => x"00000000", 28724 => x"00000000",
    28725 => x"00000000", 28726 => x"00000000", 28727 => x"00000000",
    28728 => x"00000000", 28729 => x"00000000", 28730 => x"00000000",
    28731 => x"00000000", 28732 => x"00000000", 28733 => x"00000000",
    28734 => x"00000000", 28735 => x"00000000", 28736 => x"00000000",
    28737 => x"00000000", 28738 => x"00000000", 28739 => x"00000000",
    28740 => x"00000000", 28741 => x"00000000", 28742 => x"00000000",
    28743 => x"00000000", 28744 => x"00000000", 28745 => x"00000000",
    28746 => x"00000000", 28747 => x"00000000", 28748 => x"00000000",
    28749 => x"00000000", 28750 => x"00000000", 28751 => x"00000000",
    28752 => x"00000000", 28753 => x"00000000", 28754 => x"00000000",
    28755 => x"00000000", 28756 => x"00000000", 28757 => x"00000000",
    28758 => x"00000000", 28759 => x"00000000", 28760 => x"00000000",
    28761 => x"00000000", 28762 => x"00000000", 28763 => x"00000000",
    28764 => x"00000000", 28765 => x"00000000", 28766 => x"00000000",
    28767 => x"00000000", 28768 => x"00000000", 28769 => x"00000000",
    28770 => x"00000000", 28771 => x"00000000", 28772 => x"00000000",
    28773 => x"00000000", 28774 => x"00000000", 28775 => x"00000000",
    28776 => x"00000000", 28777 => x"00000000", 28778 => x"00000000",
    28779 => x"00000000", 28780 => x"00000000", 28781 => x"00000000",
    28782 => x"00000000", 28783 => x"00000000", 28784 => x"00000000",
    28785 => x"00000000", 28786 => x"00000000", 28787 => x"00000000",
    28788 => x"00000000", 28789 => x"00000000", 28790 => x"00000000",
    28791 => x"00000000", 28792 => x"00000000", 28793 => x"00000000",
    28794 => x"00000000", 28795 => x"00000000", 28796 => x"00000000",
    28797 => x"00000000", 28798 => x"00000000", 28799 => x"00000000",
    28800 => x"00000000", 28801 => x"00000000", 28802 => x"00000000",
    28803 => x"00000000", 28804 => x"00000000", 28805 => x"00000000",
    28806 => x"00000000", 28807 => x"00000000", 28808 => x"00000000",
    28809 => x"00000000", 28810 => x"00000000", 28811 => x"00000000",
    28812 => x"00000000", 28813 => x"00000000", 28814 => x"00000000",
    28815 => x"00000000", 28816 => x"00000000", 28817 => x"00000000",
    28818 => x"00000000", 28819 => x"00000000", 28820 => x"00000000",
    28821 => x"00000000", 28822 => x"00000000", 28823 => x"00000000",
    28824 => x"00000000", 28825 => x"00000000", 28826 => x"00000000",
    28827 => x"00000000", 28828 => x"00000000", 28829 => x"00000000",
    28830 => x"00000000", 28831 => x"00000000", 28832 => x"00000000",
    28833 => x"00000000", 28834 => x"00000000", 28835 => x"00000000",
    28836 => x"00000000", 28837 => x"00000000", 28838 => x"00000000",
    28839 => x"00000000", 28840 => x"00000000", 28841 => x"00000000",
    28842 => x"00000000", 28843 => x"00000000", 28844 => x"00000000",
    28845 => x"00000000", 28846 => x"00000000", 28847 => x"00000000",
    28848 => x"00000000", 28849 => x"00000000", 28850 => x"00000000",
    28851 => x"00000000", 28852 => x"00000000", 28853 => x"00000000",
    28854 => x"00000000", 28855 => x"00000000", 28856 => x"00000000",
    28857 => x"00000000", 28858 => x"00000000", 28859 => x"00000000",
    28860 => x"00000000", 28861 => x"00000000", 28862 => x"00000000",
    28863 => x"00000000", 28864 => x"00000000", 28865 => x"00000000",
    28866 => x"00000000", 28867 => x"00000000", 28868 => x"00000000",
    28869 => x"00000000", 28870 => x"00000000", 28871 => x"00000000",
    28872 => x"00000000", 28873 => x"00000000", 28874 => x"00000000",
    28875 => x"00000000", 28876 => x"00000000", 28877 => x"00000000",
    28878 => x"00000000", 28879 => x"00000000", 28880 => x"00000000",
    28881 => x"00000000", 28882 => x"00000000", 28883 => x"00000000",
    28884 => x"00000000", 28885 => x"00000000", 28886 => x"00000000",
    28887 => x"00000000", 28888 => x"00000000", 28889 => x"00000000",
    28890 => x"00000000", 28891 => x"00000000", 28892 => x"00000000",
    28893 => x"00000000", 28894 => x"00000000", 28895 => x"00000000",
    28896 => x"00000000", 28897 => x"00000000", 28898 => x"00000000",
    28899 => x"00000000", 28900 => x"00000000", 28901 => x"00000000",
    28902 => x"00000000", 28903 => x"00000000", 28904 => x"00000000",
    28905 => x"00000000", 28906 => x"00000000", 28907 => x"00000000",
    28908 => x"00000000", 28909 => x"00000000", 28910 => x"00000000",
    28911 => x"00000000", 28912 => x"00000000", 28913 => x"00000000",
    28914 => x"00000000", 28915 => x"00000000", 28916 => x"00000000",
    28917 => x"00000000", 28918 => x"00000000", 28919 => x"00000000",
    28920 => x"00000000", 28921 => x"00000000", 28922 => x"00000000",
    28923 => x"00000000", 28924 => x"00000000", 28925 => x"00000000",
    28926 => x"00000000", 28927 => x"00000000", 28928 => x"00000000",
    28929 => x"00000000", 28930 => x"00000000", 28931 => x"00000000",
    28932 => x"00000000", 28933 => x"00000000", 28934 => x"00000000",
    28935 => x"00000000", 28936 => x"00000000", 28937 => x"00000000",
    28938 => x"00000000", 28939 => x"00000000", 28940 => x"00000000",
    28941 => x"00000000", 28942 => x"00000000", 28943 => x"00000000",
    28944 => x"00000000", 28945 => x"00000000", 28946 => x"00000000",
    28947 => x"00000000", 28948 => x"00000000", 28949 => x"00000000",
    28950 => x"00000000", 28951 => x"00000000", 28952 => x"00000000",
    28953 => x"00000000", 28954 => x"00000000", 28955 => x"00000000",
    28956 => x"00000000", 28957 => x"00000000", 28958 => x"00000000",
    28959 => x"00000000", 28960 => x"00000000", 28961 => x"00000000",
    28962 => x"00000000", 28963 => x"00000000", 28964 => x"00000000",
    28965 => x"00000000", 28966 => x"00000000", 28967 => x"00000000",
    28968 => x"00000000", 28969 => x"00000000", 28970 => x"00000000",
    28971 => x"00000000", 28972 => x"00000000", 28973 => x"00000000",
    28974 => x"00000000", 28975 => x"00000000", 28976 => x"00000000",
    28977 => x"00000000", 28978 => x"00000000", 28979 => x"00000000",
    28980 => x"00000000", 28981 => x"00000000", 28982 => x"00000000",
    28983 => x"00000000", 28984 => x"00000000", 28985 => x"00000000",
    28986 => x"00000000", 28987 => x"00000000", 28988 => x"00000000",
    28989 => x"00000000", 28990 => x"00000000", 28991 => x"00000000",
    28992 => x"00000000", 28993 => x"00000000", 28994 => x"00000000",
    28995 => x"00000000", 28996 => x"00000000", 28997 => x"00000000",
    28998 => x"00000000", 28999 => x"00000000", 29000 => x"00000000",
    29001 => x"00000000", 29002 => x"00000000", 29003 => x"00000000",
    29004 => x"00000000", 29005 => x"00000000", 29006 => x"00000000",
    29007 => x"00000000", 29008 => x"00000000", 29009 => x"00000000",
    29010 => x"00000000", 29011 => x"00000000", 29012 => x"00000000",
    29013 => x"00000000", 29014 => x"00000000", 29015 => x"00000000",
    29016 => x"00000000", 29017 => x"00000000", 29018 => x"00000000",
    29019 => x"00000000", 29020 => x"00000000", 29021 => x"00000000",
    29022 => x"00000000", 29023 => x"00000000", 29024 => x"00000000",
    29025 => x"00000000", 29026 => x"00000000", 29027 => x"00000000",
    29028 => x"00000000", 29029 => x"00000000", 29030 => x"00000000",
    29031 => x"00000000", 29032 => x"00000000", 29033 => x"00000000",
    29034 => x"00000000", 29035 => x"00000000", 29036 => x"00000000",
    29037 => x"00000000", 29038 => x"00000000", 29039 => x"00000000",
    29040 => x"00000000", 29041 => x"00000000", 29042 => x"00000000",
    29043 => x"00000000", 29044 => x"00000000", 29045 => x"00000000",
    29046 => x"00000000", 29047 => x"00000000", 29048 => x"00000000",
    29049 => x"00000000", 29050 => x"00000000", 29051 => x"00000000",
    29052 => x"00000000", 29053 => x"00000000", 29054 => x"00000000",
    29055 => x"00000000", 29056 => x"00000000", 29057 => x"00000000",
    29058 => x"00000000", 29059 => x"00000000", 29060 => x"00000000",
    29061 => x"00000000", 29062 => x"00000000", 29063 => x"00000000",
    29064 => x"00000000", 29065 => x"00000000", 29066 => x"00000000",
    29067 => x"00000000", 29068 => x"00000000", 29069 => x"00000000",
    29070 => x"00000000", 29071 => x"00000000", 29072 => x"00000000",
    29073 => x"00000000", 29074 => x"00000000", 29075 => x"00000000",
    29076 => x"00000000", 29077 => x"00000000", 29078 => x"00000000",
    29079 => x"00000000", 29080 => x"00000000", 29081 => x"00000000",
    29082 => x"00000000", 29083 => x"00000000", 29084 => x"00000000",
    29085 => x"00000000", 29086 => x"00000000", 29087 => x"00000000",
    29088 => x"00000000", 29089 => x"00000000", 29090 => x"00000000",
    29091 => x"00000000", 29092 => x"00000000", 29093 => x"00000000",
    29094 => x"00000000", 29095 => x"00000000", 29096 => x"00000000",
    29097 => x"00000000", 29098 => x"00000000", 29099 => x"00000000",
    29100 => x"00000000", 29101 => x"00000000", 29102 => x"00000000",
    29103 => x"00000000", 29104 => x"00000000", 29105 => x"00000000",
    29106 => x"00000000", 29107 => x"00000000", 29108 => x"00000000",
    29109 => x"00000000", 29110 => x"00000000", 29111 => x"00000000",
    29112 => x"00000000", 29113 => x"00000000", 29114 => x"00000000",
    29115 => x"00000000", 29116 => x"00000000", 29117 => x"00000000",
    29118 => x"00000000", 29119 => x"00000000", 29120 => x"00000000",
    29121 => x"00000000", 29122 => x"00000000", 29123 => x"00000000",
    29124 => x"00000000", 29125 => x"00000000", 29126 => x"00000000",
    29127 => x"00000000", 29128 => x"00000000", 29129 => x"00000000",
    29130 => x"00000000", 29131 => x"00000000", 29132 => x"00000000",
    29133 => x"00000000", 29134 => x"00000000", 29135 => x"00000000",
    29136 => x"00000000", 29137 => x"00000000", 29138 => x"00000000",
    29139 => x"00000000", 29140 => x"00000000", 29141 => x"00000000",
    29142 => x"00000000", 29143 => x"00000000", 29144 => x"00000000",
    29145 => x"00000000", 29146 => x"00000000", 29147 => x"00000000",
    29148 => x"00000000", 29149 => x"00000000", 29150 => x"00000000",
    29151 => x"00000000", 29152 => x"00000000", 29153 => x"00000000",
    29154 => x"00000000", 29155 => x"00000000", 29156 => x"00000000",
    29157 => x"00000000", 29158 => x"00000000", 29159 => x"00000000",
    29160 => x"00000000", 29161 => x"00000000", 29162 => x"00000000",
    29163 => x"00000000", 29164 => x"00000000", 29165 => x"00000000",
    29166 => x"00000000", 29167 => x"00000000", 29168 => x"00000000",
    29169 => x"00000000", 29170 => x"00000000", 29171 => x"00000000",
    29172 => x"00000000", 29173 => x"00000000", 29174 => x"00000000",
    29175 => x"00000000", 29176 => x"00000000", 29177 => x"00000000",
    29178 => x"00000000", 29179 => x"00000000", 29180 => x"00000000",
    29181 => x"00000000", 29182 => x"00000000", 29183 => x"00000000",
    29184 => x"00000000", 29185 => x"00000000", 29186 => x"00000000",
    29187 => x"00000000", 29188 => x"00000000", 29189 => x"00000000",
    29190 => x"00000000", 29191 => x"00000000", 29192 => x"00000000",
    29193 => x"00000000", 29194 => x"00000000", 29195 => x"00000000",
    29196 => x"00000000", 29197 => x"00000000", 29198 => x"00000000",
    29199 => x"00000000", 29200 => x"00000000", 29201 => x"00000000",
    29202 => x"00000000", 29203 => x"00000000", 29204 => x"00000000",
    29205 => x"00000000", 29206 => x"00000000", 29207 => x"00000000",
    29208 => x"00000000", 29209 => x"00000000", 29210 => x"00000000",
    29211 => x"00000000", 29212 => x"00000000", 29213 => x"00000000",
    29214 => x"00000000", 29215 => x"00000000", 29216 => x"00000000",
    29217 => x"00000000", 29218 => x"00000000", 29219 => x"00000000",
    29220 => x"00000000", 29221 => x"00000000", 29222 => x"00000000",
    29223 => x"00000000", 29224 => x"00000000", 29225 => x"00000000",
    29226 => x"00000000", 29227 => x"00000000", 29228 => x"00000000",
    29229 => x"00000000", 29230 => x"00000000", 29231 => x"00000000",
    29232 => x"00000000", 29233 => x"00000000", 29234 => x"00000000",
    29235 => x"00000000", 29236 => x"00000000", 29237 => x"00000000",
    29238 => x"00000000", 29239 => x"00000000", 29240 => x"00000000",
    29241 => x"00000000", 29242 => x"00000000", 29243 => x"00000000",
    29244 => x"00000000", 29245 => x"00000000", 29246 => x"00000000",
    29247 => x"00000000", 29248 => x"00000000", 29249 => x"00000000",
    29250 => x"00000000", 29251 => x"00000000", 29252 => x"00000000",
    29253 => x"00000000", 29254 => x"00000000", 29255 => x"00000000",
    29256 => x"00000000", 29257 => x"00000000", 29258 => x"00000000",
    29259 => x"00000000", 29260 => x"00000000", 29261 => x"00000000",
    29262 => x"00000000", 29263 => x"00000000", 29264 => x"00000000",
    29265 => x"00000000", 29266 => x"00000000", 29267 => x"00000000",
    29268 => x"00000000", 29269 => x"00000000", 29270 => x"00000000",
    29271 => x"00000000", 29272 => x"00000000", 29273 => x"00000000",
    29274 => x"00000000", 29275 => x"00000000", 29276 => x"00000000",
    29277 => x"00000000", 29278 => x"00000000", 29279 => x"00000000",
    29280 => x"00000000", 29281 => x"00000000", 29282 => x"00000000",
    29283 => x"00000000", 29284 => x"00000000", 29285 => x"00000000",
    29286 => x"00000000", 29287 => x"00000000", 29288 => x"00000000",
    29289 => x"00000000", 29290 => x"00000000", 29291 => x"00000000",
    29292 => x"00000000", 29293 => x"00000000", 29294 => x"00000000",
    29295 => x"00000000", 29296 => x"00000000", 29297 => x"00000000",
    29298 => x"00000000", 29299 => x"00000000", 29300 => x"00000000",
    29301 => x"00000000", 29302 => x"00000000", 29303 => x"00000000",
    29304 => x"00000000", 29305 => x"00000000", 29306 => x"00000000",
    29307 => x"00000000", 29308 => x"00000000", 29309 => x"00000000",
    29310 => x"00000000", 29311 => x"00000000", 29312 => x"00000000",
    29313 => x"00000000", 29314 => x"00000000", 29315 => x"00000000",
    29316 => x"00000000", 29317 => x"00000000", 29318 => x"00000000",
    29319 => x"00000000", 29320 => x"00000000", 29321 => x"00000000",
    29322 => x"00000000", 29323 => x"00000000", 29324 => x"00000000",
    29325 => x"00000000", 29326 => x"00000000", 29327 => x"00000000",
    29328 => x"00000000", 29329 => x"00000000", 29330 => x"00000000",
    29331 => x"00000000", 29332 => x"00000000", 29333 => x"00000000",
    29334 => x"00000000", 29335 => x"00000000", 29336 => x"00000000",
    29337 => x"00000000", 29338 => x"00000000", 29339 => x"00000000",
    29340 => x"00000000", 29341 => x"00000000", 29342 => x"00000000",
    29343 => x"00000000", 29344 => x"00000000", 29345 => x"00000000",
    29346 => x"00000000", 29347 => x"00000000", 29348 => x"00000000",
    29349 => x"00000000", 29350 => x"00000000", 29351 => x"00000000",
    29352 => x"00000000", 29353 => x"00000000", 29354 => x"00000000",
    29355 => x"00000000", 29356 => x"00000000", 29357 => x"00000000",
    29358 => x"00000000", 29359 => x"00000000", 29360 => x"00000000",
    29361 => x"00000000", 29362 => x"00000000", 29363 => x"00000000",
    29364 => x"00000000", 29365 => x"00000000", 29366 => x"00000000",
    29367 => x"00000000", 29368 => x"00000000", 29369 => x"00000000",
    29370 => x"00000000", 29371 => x"00000000", 29372 => x"00000000",
    29373 => x"00000000", 29374 => x"00000000", 29375 => x"00000000",
    29376 => x"00000000", 29377 => x"00000000", 29378 => x"00000000",
    29379 => x"00000000", 29380 => x"00000000", 29381 => x"00000000",
    29382 => x"00000000", 29383 => x"00000000", 29384 => x"00000000",
    29385 => x"00000000", 29386 => x"00000000", 29387 => x"00000000",
    29388 => x"00000000", 29389 => x"00000000", 29390 => x"00000000",
    29391 => x"00000000", 29392 => x"00000000", 29393 => x"00000000",
    29394 => x"00000000", 29395 => x"00000000", 29396 => x"00000000",
    29397 => x"00000000", 29398 => x"00000000", 29399 => x"00000000",
    29400 => x"00000000", 29401 => x"00000000", 29402 => x"00000000",
    29403 => x"00000000", 29404 => x"00000000", 29405 => x"00000000",
    29406 => x"00000000", 29407 => x"00000000", 29408 => x"00000000",
    29409 => x"00000000", 29410 => x"00000000", 29411 => x"00000000",
    29412 => x"00000000", 29413 => x"00000000", 29414 => x"00000000",
    29415 => x"00000000", 29416 => x"00000000", 29417 => x"00000000",
    29418 => x"00000000", 29419 => x"00000000", 29420 => x"00000000",
    29421 => x"00000000", 29422 => x"00000000", 29423 => x"00000000",
    29424 => x"00000000", 29425 => x"00000000", 29426 => x"00000000",
    29427 => x"00000000", 29428 => x"00000000", 29429 => x"00000000",
    29430 => x"00000000", 29431 => x"00000000", 29432 => x"00000000",
    29433 => x"00000000", 29434 => x"00000000", 29435 => x"00000000",
    29436 => x"00000000", 29437 => x"00000000", 29438 => x"00000000",
    29439 => x"00000000", 29440 => x"00000000", 29441 => x"00000000",
    29442 => x"00000000", 29443 => x"00000000", 29444 => x"00000000",
    29445 => x"00000000", 29446 => x"00000000", 29447 => x"00000000",
    29448 => x"00000000", 29449 => x"00000000", 29450 => x"00000000",
    29451 => x"00000000", 29452 => x"00000000", 29453 => x"00000000",
    29454 => x"00000000", 29455 => x"00000000", 29456 => x"00000000",
    29457 => x"00000000", 29458 => x"00000000", 29459 => x"00000000",
    29460 => x"00000000", 29461 => x"00000000", 29462 => x"00000000",
    29463 => x"00000000", 29464 => x"00000000", 29465 => x"00000000",
    29466 => x"00000000", 29467 => x"00000000", 29468 => x"00000000",
    29469 => x"00000000", 29470 => x"00000000", 29471 => x"00000000",
    29472 => x"00000000", 29473 => x"00000000", 29474 => x"00000000",
    29475 => x"00000000", 29476 => x"00000000", 29477 => x"00000000",
    29478 => x"00000000", 29479 => x"00000000", 29480 => x"00000000",
    29481 => x"00000000", 29482 => x"00000000", 29483 => x"00000000",
    29484 => x"00000000", 29485 => x"00000000", 29486 => x"00000000",
    29487 => x"00000000", 29488 => x"00000000", 29489 => x"00000000",
    29490 => x"00000000", 29491 => x"00000000", 29492 => x"00000000",
    29493 => x"00000000", 29494 => x"00000000", 29495 => x"00000000",
    29496 => x"00000000", 29497 => x"00000000", 29498 => x"00000000",
    29499 => x"00000000", 29500 => x"00000000", 29501 => x"00000000",
    29502 => x"00000000", 29503 => x"00000000", 29504 => x"00000000",
    29505 => x"00000000", 29506 => x"00000000", 29507 => x"00000000",
    29508 => x"00000000", 29509 => x"00000000", 29510 => x"00000000",
    29511 => x"00000000", 29512 => x"00000000", 29513 => x"00000000",
    29514 => x"00000000", 29515 => x"00000000", 29516 => x"00000000",
    29517 => x"00000000", 29518 => x"00000000", 29519 => x"00000000",
    29520 => x"00000000", 29521 => x"00000000", 29522 => x"00000000",
    29523 => x"00000000", 29524 => x"00000000", 29525 => x"00000000",
    29526 => x"00000000", 29527 => x"00000000", 29528 => x"00000000",
    29529 => x"00000000", 29530 => x"00000000", 29531 => x"00000000",
    29532 => x"00000000", 29533 => x"00000000", 29534 => x"00000000",
    29535 => x"00000000", 29536 => x"00000000", 29537 => x"00000000",
    29538 => x"00000000", 29539 => x"00000000", 29540 => x"00000000",
    29541 => x"00000000", 29542 => x"00000000", 29543 => x"00000000",
    29544 => x"00000000", 29545 => x"00000000", 29546 => x"00000000",
    29547 => x"00000000", 29548 => x"00000000", 29549 => x"00000000",
    29550 => x"00000000", 29551 => x"00000000", 29552 => x"00000000",
    29553 => x"00000000", 29554 => x"00000000", 29555 => x"00000000",
    29556 => x"00000000", 29557 => x"00000000", 29558 => x"00000000",
    29559 => x"00000000", 29560 => x"00000000", 29561 => x"00000000",
    29562 => x"00000000", 29563 => x"00000000", 29564 => x"00000000",
    29565 => x"00000000", 29566 => x"00000000", 29567 => x"00000000",
    29568 => x"00000000", 29569 => x"00000000", 29570 => x"00000000",
    29571 => x"00000000", 29572 => x"00000000", 29573 => x"00000000",
    29574 => x"00000000", 29575 => x"00000000", 29576 => x"00000000",
    29577 => x"00000000", 29578 => x"00000000", 29579 => x"00000000",
    29580 => x"00000000", 29581 => x"00000000", 29582 => x"00000000",
    29583 => x"00000000", 29584 => x"00000000", 29585 => x"00000000",
    29586 => x"00000000", 29587 => x"00000000", 29588 => x"00000000",
    29589 => x"00000000", 29590 => x"00000000", 29591 => x"00000000",
    29592 => x"00000000", 29593 => x"00000000", 29594 => x"00000000",
    29595 => x"00000000", 29596 => x"00000000", 29597 => x"00000000",
    29598 => x"00000000", 29599 => x"00000000", 29600 => x"00000000",
    29601 => x"00000000", 29602 => x"00000000", 29603 => x"00000000",
    29604 => x"00000000", 29605 => x"00000000", 29606 => x"00000000",
    29607 => x"00000000", 29608 => x"00000000", 29609 => x"00000000",
    29610 => x"00000000", 29611 => x"00000000", 29612 => x"00000000",
    29613 => x"00000000", 29614 => x"00000000", 29615 => x"00000000",
    29616 => x"00000000", 29617 => x"00000000", 29618 => x"00000000",
    29619 => x"00000000", 29620 => x"00000000", 29621 => x"00000000",
    29622 => x"00000000", 29623 => x"00000000", 29624 => x"00000000",
    29625 => x"00000000", 29626 => x"00000000", 29627 => x"00000000",
    29628 => x"00000000", 29629 => x"00000000", 29630 => x"00000000",
    29631 => x"00000000", 29632 => x"00000000", 29633 => x"00000000",
    29634 => x"00000000", 29635 => x"00000000", 29636 => x"00000000",
    29637 => x"00000000", 29638 => x"00000000", 29639 => x"00000000",
    29640 => x"00000000", 29641 => x"00000000", 29642 => x"00000000",
    29643 => x"00000000", 29644 => x"00000000", 29645 => x"00000000",
    29646 => x"00000000", 29647 => x"00000000", 29648 => x"00000000",
    29649 => x"00000000", 29650 => x"00000000", 29651 => x"00000000",
    29652 => x"00000000", 29653 => x"00000000", 29654 => x"00000000",
    29655 => x"00000000", 29656 => x"00000000", 29657 => x"00000000",
    29658 => x"00000000", 29659 => x"00000000", 29660 => x"00000000",
    29661 => x"00000000", 29662 => x"00000000", 29663 => x"00000000",
    29664 => x"00000000", 29665 => x"00000000", 29666 => x"00000000",
    29667 => x"00000000", 29668 => x"00000000", 29669 => x"00000000",
    29670 => x"00000000", 29671 => x"00000000", 29672 => x"00000000",
    29673 => x"00000000", 29674 => x"00000000", 29675 => x"00000000",
    29676 => x"00000000", 29677 => x"00000000", 29678 => x"00000000",
    29679 => x"00000000", 29680 => x"00000000", 29681 => x"00000000",
    29682 => x"00000000", 29683 => x"00000000", 29684 => x"00000000",
    29685 => x"00000000", 29686 => x"00000000", 29687 => x"00000000",
    29688 => x"00000000", 29689 => x"00000000", 29690 => x"00000000",
    29691 => x"00000000", 29692 => x"00000000", 29693 => x"00000000",
    29694 => x"00000000", 29695 => x"00000000", 29696 => x"00000000",
    29697 => x"00000000", 29698 => x"00000000", 29699 => x"00000000",
    29700 => x"00000000", 29701 => x"00000000", 29702 => x"00000000",
    29703 => x"00000000", 29704 => x"00000000", 29705 => x"00000000",
    29706 => x"00000000", 29707 => x"00000000", 29708 => x"00000000",
    29709 => x"00000000", 29710 => x"00000000", 29711 => x"00000000",
    29712 => x"00000000", 29713 => x"00000000", 29714 => x"00000000",
    29715 => x"00000000", 29716 => x"00000000", 29717 => x"00000000",
    29718 => x"00000000", 29719 => x"00000000", 29720 => x"00000000",
    29721 => x"00000000", 29722 => x"00000000", 29723 => x"00000000",
    29724 => x"00000000", 29725 => x"00000000", 29726 => x"00000000",
    29727 => x"00000000", 29728 => x"00000000", 29729 => x"00000000",
    29730 => x"00000000", 29731 => x"00000000", 29732 => x"00000000",
    29733 => x"00000000", 29734 => x"00000000", 29735 => x"00000000",
    29736 => x"00000000", 29737 => x"00000000", 29738 => x"00000000",
    29739 => x"00000000", 29740 => x"00000000", 29741 => x"00000000",
    29742 => x"00000000", 29743 => x"00000000", 29744 => x"00000000",
    29745 => x"00000000", 29746 => x"00000000", 29747 => x"00000000",
    29748 => x"00000000", 29749 => x"00000000", 29750 => x"00000000",
    29751 => x"00000000", 29752 => x"00000000", 29753 => x"00000000",
    29754 => x"00000000", 29755 => x"00000000", 29756 => x"00000000",
    29757 => x"00000000", 29758 => x"00000000", 29759 => x"00000000",
    29760 => x"00000000", 29761 => x"00000000", 29762 => x"00000000",
    29763 => x"00000000", 29764 => x"00000000", 29765 => x"00000000",
    29766 => x"00000000", 29767 => x"00000000", 29768 => x"00000000",
    29769 => x"00000000", 29770 => x"00000000", 29771 => x"00000000",
    29772 => x"00000000", 29773 => x"00000000", 29774 => x"00000000",
    29775 => x"00000000", 29776 => x"00000000", 29777 => x"00000000",
    29778 => x"00000000", 29779 => x"00000000", 29780 => x"00000000",
    29781 => x"00000000", 29782 => x"00000000", 29783 => x"00000000",
    29784 => x"00000000", 29785 => x"00000000", 29786 => x"00000000",
    29787 => x"00000000", 29788 => x"00000000", 29789 => x"00000000",
    29790 => x"00000000", 29791 => x"00000000", 29792 => x"00000000",
    29793 => x"00000000", 29794 => x"00000000", 29795 => x"00000000",
    29796 => x"00000000", 29797 => x"00000000", 29798 => x"00000000",
    29799 => x"00000000", 29800 => x"00000000", 29801 => x"00000000",
    29802 => x"00000000", 29803 => x"00000000", 29804 => x"00000000",
    29805 => x"00000000", 29806 => x"00000000", 29807 => x"00000000",
    29808 => x"00000000", 29809 => x"00000000", 29810 => x"00000000",
    29811 => x"00000000", 29812 => x"00000000", 29813 => x"00000000",
    29814 => x"00000000", 29815 => x"00000000", 29816 => x"00000000",
    29817 => x"00000000", 29818 => x"00000000", 29819 => x"00000000",
    29820 => x"00000000", 29821 => x"00000000", 29822 => x"00000000",
    29823 => x"00000000", 29824 => x"00000000", 29825 => x"00000000",
    29826 => x"00000000", 29827 => x"00000000", 29828 => x"00000000",
    29829 => x"00000000", 29830 => x"00000000", 29831 => x"00000000",
    29832 => x"00000000", 29833 => x"00000000", 29834 => x"00000000",
    29835 => x"00000000", 29836 => x"00000000", 29837 => x"00000000",
    29838 => x"00000000", 29839 => x"00000000", 29840 => x"00000000",
    29841 => x"00000000", 29842 => x"00000000", 29843 => x"00000000",
    29844 => x"00000000", 29845 => x"00000000", 29846 => x"00000000",
    29847 => x"00000000", 29848 => x"00000000", 29849 => x"00000000",
    29850 => x"00000000", 29851 => x"00000000", 29852 => x"00000000",
    29853 => x"00000000", 29854 => x"00000000", 29855 => x"00000000",
    29856 => x"00000000", 29857 => x"00000000", 29858 => x"00000000",
    29859 => x"00000000", 29860 => x"00000000", 29861 => x"00000000",
    29862 => x"00000000", 29863 => x"00000000", 29864 => x"00000000",
    29865 => x"00000000", 29866 => x"00000000", 29867 => x"00000000",
    29868 => x"00000000", 29869 => x"00000000", 29870 => x"00000000",
    29871 => x"00000000", 29872 => x"00000000", 29873 => x"00000000",
    29874 => x"00000000", 29875 => x"00000000", 29876 => x"00000000",
    29877 => x"00000000", 29878 => x"00000000", 29879 => x"00000000",
    29880 => x"00000000", 29881 => x"00000000", 29882 => x"00000000",
    29883 => x"00000000", 29884 => x"00000000", 29885 => x"00000000",
    29886 => x"00000000", 29887 => x"00000000", 29888 => x"00000000",
    29889 => x"00000000", 29890 => x"00000000", 29891 => x"00000000",
    29892 => x"00000000", 29893 => x"00000000", 29894 => x"00000000",
    29895 => x"00000000", 29896 => x"00000000", 29897 => x"00000000",
    29898 => x"00000000", 29899 => x"00000000", 29900 => x"00000000",
    29901 => x"00000000", 29902 => x"00000000", 29903 => x"00000000",
    29904 => x"00000000", 29905 => x"00000000", 29906 => x"00000000",
    29907 => x"00000000", 29908 => x"00000000", 29909 => x"00000000",
    29910 => x"00000000", 29911 => x"00000000", 29912 => x"00000000",
    29913 => x"00000000", 29914 => x"00000000", 29915 => x"00000000",
    29916 => x"00000000", 29917 => x"00000000", 29918 => x"00000000",
    29919 => x"00000000", 29920 => x"00000000", 29921 => x"00000000",
    29922 => x"00000000", 29923 => x"00000000", 29924 => x"00000000",
    29925 => x"00000000", 29926 => x"00000000", 29927 => x"00000000",
    29928 => x"00000000", 29929 => x"00000000", 29930 => x"00000000",
    29931 => x"00000000", 29932 => x"00000000", 29933 => x"00000000",
    29934 => x"00000000", 29935 => x"00000000", 29936 => x"00000000",
    29937 => x"00000000", 29938 => x"00000000", 29939 => x"00000000",
    29940 => x"00000000", 29941 => x"00000000", 29942 => x"00000000",
    29943 => x"00000000", 29944 => x"00000000", 29945 => x"00000000",
    29946 => x"00000000", 29947 => x"00000000", 29948 => x"00000000",
    29949 => x"00000000", 29950 => x"00000000", 29951 => x"00000000",
    29952 => x"00000000", 29953 => x"00000000", 29954 => x"00000000",
    29955 => x"00000000", 29956 => x"00000000", 29957 => x"00000000",
    29958 => x"00000000", 29959 => x"00000000", 29960 => x"00000000",
    29961 => x"00000000", 29962 => x"00000000", 29963 => x"00000000",
    29964 => x"00000000", 29965 => x"00000000", 29966 => x"00000000",
    29967 => x"00000000", 29968 => x"00000000", 29969 => x"00000000",
    29970 => x"00000000", 29971 => x"00000000", 29972 => x"00000000",
    29973 => x"00000000", 29974 => x"00000000", 29975 => x"00000000",
    29976 => x"00000000", 29977 => x"00000000", 29978 => x"00000000",
    29979 => x"00000000", 29980 => x"00000000", 29981 => x"00000000",
    29982 => x"00000000", 29983 => x"00000000", 29984 => x"00000000",
    29985 => x"00000000", 29986 => x"00000000", 29987 => x"00000000",
    29988 => x"00000000", 29989 => x"00000000", 29990 => x"00000000",
    29991 => x"00000000", 29992 => x"00000000", 29993 => x"00000000",
    29994 => x"00000000", 29995 => x"00000000", 29996 => x"00000000",
    29997 => x"00000000", 29998 => x"00000000", 29999 => x"00000000",
    30000 => x"00000000", 30001 => x"00000000", 30002 => x"00000000",
    30003 => x"00000000", 30004 => x"00000000", 30005 => x"00000000",
    30006 => x"00000000", 30007 => x"00000000", 30008 => x"00000000",
    30009 => x"00000000", 30010 => x"00000000", 30011 => x"00000000",
    30012 => x"00000000", 30013 => x"00000000", 30014 => x"00000000",
    30015 => x"00000000", 30016 => x"00000000", 30017 => x"00000000",
    30018 => x"00000000", 30019 => x"00000000", 30020 => x"00000000",
    30021 => x"00000000", 30022 => x"00000000", 30023 => x"00000000",
    30024 => x"00000000", 30025 => x"00000000", 30026 => x"00000000",
    30027 => x"00000000", 30028 => x"00000000", 30029 => x"00000000",
    30030 => x"00000000", 30031 => x"00000000", 30032 => x"00000000",
    30033 => x"00000000", 30034 => x"00000000", 30035 => x"00000000",
    30036 => x"00000000", 30037 => x"00000000", 30038 => x"00000000",
    30039 => x"00000000", 30040 => x"00000000", 30041 => x"00000000",
    30042 => x"00000000", 30043 => x"00000000", 30044 => x"00000000",
    30045 => x"00000000", 30046 => x"00000000", 30047 => x"00000000",
    30048 => x"00000000", 30049 => x"00000000", 30050 => x"00000000",
    30051 => x"00000000", 30052 => x"00000000", 30053 => x"00000000",
    30054 => x"00000000", 30055 => x"00000000", 30056 => x"00000000",
    30057 => x"00000000", 30058 => x"00000000", 30059 => x"00000000",
    30060 => x"00000000", 30061 => x"00000000", 30062 => x"00000000",
    30063 => x"00000000", 30064 => x"00000000", 30065 => x"00000000",
    30066 => x"00000000", 30067 => x"00000000", 30068 => x"00000000",
    30069 => x"00000000", 30070 => x"00000000", 30071 => x"00000000",
    30072 => x"00000000", 30073 => x"00000000", 30074 => x"00000000",
    30075 => x"00000000", 30076 => x"00000000", 30077 => x"00000000",
    30078 => x"00000000", 30079 => x"00000000", 30080 => x"00000000",
    30081 => x"00000000", 30082 => x"00000000", 30083 => x"00000000",
    30084 => x"00000000", 30085 => x"00000000", 30086 => x"00000000",
    30087 => x"00000000", 30088 => x"00000000", 30089 => x"00000000",
    30090 => x"00000000", 30091 => x"00000000", 30092 => x"00000000",
    30093 => x"00000000", 30094 => x"00000000", 30095 => x"00000000",
    30096 => x"00000000", 30097 => x"00000000", 30098 => x"00000000",
    30099 => x"00000000", 30100 => x"00000000", 30101 => x"00000000",
    30102 => x"00000000", 30103 => x"00000000", 30104 => x"00000000",
    30105 => x"00000000", 30106 => x"00000000", 30107 => x"00000000",
    30108 => x"00000000", 30109 => x"00000000", 30110 => x"00000000",
    30111 => x"00000000", 30112 => x"00000000", 30113 => x"00000000",
    30114 => x"00000000", 30115 => x"00000000", 30116 => x"00000000",
    30117 => x"00000000", 30118 => x"00000000", 30119 => x"00000000",
    30120 => x"00000000", 30121 => x"00000000", 30122 => x"00000000",
    30123 => x"00000000", 30124 => x"00000000", 30125 => x"00000000",
    30126 => x"00000000", 30127 => x"00000000", 30128 => x"00000000",
    30129 => x"00000000", 30130 => x"00000000", 30131 => x"00000000",
    30132 => x"00000000", 30133 => x"00000000", 30134 => x"00000000",
    30135 => x"00000000", 30136 => x"00000000", 30137 => x"00000000",
    30138 => x"00000000", 30139 => x"00000000", 30140 => x"00000000",
    30141 => x"00000000", 30142 => x"00000000", 30143 => x"00000000",
    30144 => x"00000000", 30145 => x"00000000", 30146 => x"00000000",
    30147 => x"00000000", 30148 => x"00000000", 30149 => x"00000000",
    30150 => x"00000000", 30151 => x"00000000", 30152 => x"00000000",
    30153 => x"00000000", 30154 => x"00000000", 30155 => x"00000000",
    30156 => x"00000000", 30157 => x"00000000", 30158 => x"00000000",
    30159 => x"00000000", 30160 => x"00000000", 30161 => x"00000000",
    30162 => x"00000000", 30163 => x"00000000", 30164 => x"00000000",
    30165 => x"00000000", 30166 => x"00000000", 30167 => x"00000000",
    30168 => x"00000000", 30169 => x"00000000", 30170 => x"00000000",
    30171 => x"00000000", 30172 => x"00000000", 30173 => x"00000000",
    30174 => x"00000000", 30175 => x"00000000", 30176 => x"00000000",
    30177 => x"00000000", 30178 => x"00000000", 30179 => x"00000000",
    30180 => x"00000000", 30181 => x"00000000", 30182 => x"00000000",
    30183 => x"00000000", 30184 => x"00000000", 30185 => x"00000000",
    30186 => x"00000000", 30187 => x"00000000", 30188 => x"00000000",
    30189 => x"00000000", 30190 => x"00000000", 30191 => x"00000000",
    30192 => x"00000000", 30193 => x"00000000", 30194 => x"00000000",
    30195 => x"00000000", 30196 => x"00000000", 30197 => x"00000000",
    30198 => x"00000000", 30199 => x"00000000", 30200 => x"00000000",
    30201 => x"00000000", 30202 => x"00000000", 30203 => x"00000000",
    30204 => x"00000000", 30205 => x"00000000", 30206 => x"00000000",
    30207 => x"00000000", 30208 => x"00000000", 30209 => x"00000000",
    30210 => x"00000000", 30211 => x"00000000", 30212 => x"00000000",
    30213 => x"00000000", 30214 => x"00000000", 30215 => x"00000000",
    30216 => x"00000000", 30217 => x"00000000", 30218 => x"00000000",
    30219 => x"00000000", 30220 => x"00000000", 30221 => x"00000000",
    30222 => x"00000000", 30223 => x"00000000", 30224 => x"00000000",
    30225 => x"00000000", 30226 => x"00000000", 30227 => x"00000000",
    30228 => x"00000000", 30229 => x"00000000", 30230 => x"00000000",
    30231 => x"00000000", 30232 => x"00000000", 30233 => x"00000000",
    30234 => x"00000000", 30235 => x"00000000", 30236 => x"00000000",
    30237 => x"00000000", 30238 => x"00000000", 30239 => x"00000000",
    30240 => x"00000000", 30241 => x"00000000", 30242 => x"00000000",
    30243 => x"00000000", 30244 => x"00000000", 30245 => x"00000000",
    30246 => x"00000000", 30247 => x"00000000", 30248 => x"00000000",
    30249 => x"00000000", 30250 => x"00000000", 30251 => x"00000000",
    30252 => x"00000000", 30253 => x"00000000", 30254 => x"00000000",
    30255 => x"00000000", 30256 => x"00000000", 30257 => x"00000000",
    30258 => x"00000000", 30259 => x"00000000", 30260 => x"00000000",
    30261 => x"00000000", 30262 => x"00000000", 30263 => x"00000000",
    30264 => x"00000000", 30265 => x"00000000", 30266 => x"00000000",
    30267 => x"00000000", 30268 => x"00000000", 30269 => x"00000000",
    30270 => x"00000000", 30271 => x"00000000", 30272 => x"00000000",
    30273 => x"00000000", 30274 => x"00000000", 30275 => x"00000000",
    30276 => x"00000000", 30277 => x"00000000", 30278 => x"00000000",
    30279 => x"00000000", 30280 => x"00000000", 30281 => x"00000000",
    30282 => x"00000000", 30283 => x"00000000", 30284 => x"00000000",
    30285 => x"00000000", 30286 => x"00000000", 30287 => x"00000000",
    30288 => x"00000000", 30289 => x"00000000", 30290 => x"00000000",
    30291 => x"00000000", 30292 => x"00000000", 30293 => x"00000000",
    30294 => x"00000000", 30295 => x"00000000", 30296 => x"00000000",
    30297 => x"00000000", 30298 => x"00000000", 30299 => x"00000000",
    30300 => x"00000000", 30301 => x"00000000", 30302 => x"00000000",
    30303 => x"00000000", 30304 => x"00000000", 30305 => x"00000000",
    30306 => x"00000000", 30307 => x"00000000", 30308 => x"00000000",
    30309 => x"00000000", 30310 => x"00000000", 30311 => x"00000000",
    30312 => x"00000000", 30313 => x"00000000", 30314 => x"00000000",
    30315 => x"00000000", 30316 => x"00000000", 30317 => x"00000000",
    30318 => x"00000000", 30319 => x"00000000", 30320 => x"00000000",
    30321 => x"00000000", 30322 => x"00000000", 30323 => x"00000000",
    30324 => x"00000000", 30325 => x"00000000", 30326 => x"00000000",
    30327 => x"00000000", 30328 => x"00000000", 30329 => x"00000000",
    30330 => x"00000000", 30331 => x"00000000", 30332 => x"00000000",
    30333 => x"00000000", 30334 => x"00000000", 30335 => x"00000000",
    30336 => x"00000000", 30337 => x"00000000", 30338 => x"00000000",
    30339 => x"00000000", 30340 => x"00000000", 30341 => x"00000000",
    30342 => x"00000000", 30343 => x"00000000", 30344 => x"00000000",
    30345 => x"00000000", 30346 => x"00000000", 30347 => x"00000000",
    30348 => x"00000000", 30349 => x"00000000", 30350 => x"00000000",
    30351 => x"00000000", 30352 => x"00000000", 30353 => x"00000000",
    30354 => x"00000000", 30355 => x"00000000", 30356 => x"00000000",
    30357 => x"00000000", 30358 => x"00000000", 30359 => x"00000000",
    30360 => x"00000000", 30361 => x"00000000", 30362 => x"00000000",
    30363 => x"00000000", 30364 => x"00000000", 30365 => x"00000000",
    30366 => x"00000000", 30367 => x"00000000", 30368 => x"00000000",
    30369 => x"00000000", 30370 => x"00000000", 30371 => x"00000000",
    30372 => x"00000000", 30373 => x"00000000", 30374 => x"00000000",
    30375 => x"00000000", 30376 => x"00000000", 30377 => x"00000000",
    30378 => x"00000000", 30379 => x"00000000", 30380 => x"00000000",
    30381 => x"00000000", 30382 => x"00000000", 30383 => x"00000000",
    30384 => x"00000000", 30385 => x"00000000", 30386 => x"00000000",
    30387 => x"00000000", 30388 => x"00000000", 30389 => x"00000000",
    30390 => x"00000000", 30391 => x"00000000", 30392 => x"00000000",
    30393 => x"00000000", 30394 => x"00000000", 30395 => x"00000000",
    30396 => x"00000000", 30397 => x"00000000", 30398 => x"00000000",
    30399 => x"00000000", 30400 => x"00000000", 30401 => x"00000000",
    30402 => x"00000000", 30403 => x"00000000", 30404 => x"00000000",
    30405 => x"00000000", 30406 => x"00000000", 30407 => x"00000000",
    30408 => x"00000000", 30409 => x"00000000", 30410 => x"00000000",
    30411 => x"00000000", 30412 => x"00000000", 30413 => x"00000000",
    30414 => x"00000000", 30415 => x"00000000", 30416 => x"00000000",
    30417 => x"00000000", 30418 => x"00000000", 30419 => x"00000000",
    30420 => x"00000000", 30421 => x"00000000", 30422 => x"00000000",
    30423 => x"00000000", 30424 => x"00000000", 30425 => x"00000000",
    30426 => x"00000000", 30427 => x"00000000", 30428 => x"00000000",
    30429 => x"00000000", 30430 => x"00000000", 30431 => x"00000000",
    30432 => x"00000000", 30433 => x"00000000", 30434 => x"00000000",
    30435 => x"00000000", 30436 => x"00000000", 30437 => x"00000000",
    30438 => x"00000000", 30439 => x"00000000", 30440 => x"00000000",
    30441 => x"00000000", 30442 => x"00000000", 30443 => x"00000000",
    30444 => x"00000000", 30445 => x"00000000", 30446 => x"00000000",
    30447 => x"00000000", 30448 => x"00000000", 30449 => x"00000000",
    30450 => x"00000000", 30451 => x"00000000", 30452 => x"00000000",
    30453 => x"00000000", 30454 => x"00000000", 30455 => x"00000000",
    30456 => x"00000000", 30457 => x"00000000", 30458 => x"00000000",
    30459 => x"00000000", 30460 => x"00000000", 30461 => x"00000000",
    30462 => x"00000000", 30463 => x"00000000", 30464 => x"00000000",
    30465 => x"00000000", 30466 => x"00000000", 30467 => x"00000000",
    30468 => x"00000000", 30469 => x"00000000", 30470 => x"00000000",
    30471 => x"00000000", 30472 => x"00000000", 30473 => x"00000000",
    30474 => x"00000000", 30475 => x"00000000", 30476 => x"00000000",
    30477 => x"00000000", 30478 => x"00000000", 30479 => x"00000000",
    30480 => x"00000000", 30481 => x"00000000", 30482 => x"00000000",
    30483 => x"00000000", 30484 => x"00000000", 30485 => x"00000000",
    30486 => x"00000000", 30487 => x"00000000", 30488 => x"00000000",
    30489 => x"00000000", 30490 => x"00000000", 30491 => x"00000000",
    30492 => x"00000000", 30493 => x"00000000", 30494 => x"00000000",
    30495 => x"00000000", 30496 => x"00000000", 30497 => x"00000000",
    30498 => x"00000000", 30499 => x"00000000", 30500 => x"00000000",
    30501 => x"00000000", 30502 => x"00000000", 30503 => x"00000000",
    30504 => x"00000000", 30505 => x"00000000", 30506 => x"00000000",
    30507 => x"00000000", 30508 => x"00000000", 30509 => x"00000000",
    30510 => x"00000000", 30511 => x"00000000", 30512 => x"00000000",
    30513 => x"00000000", 30514 => x"00000000", 30515 => x"00000000",
    30516 => x"00000000", 30517 => x"00000000", 30518 => x"00000000",
    30519 => x"00000000", 30520 => x"00000000", 30521 => x"00000000",
    30522 => x"00000000", 30523 => x"00000000", 30524 => x"00000000",
    30525 => x"00000000", 30526 => x"00000000", 30527 => x"00000000",
    30528 => x"00000000", 30529 => x"00000000", 30530 => x"00000000",
    30531 => x"00000000", 30532 => x"00000000", 30533 => x"00000000",
    30534 => x"00000000", 30535 => x"00000000", 30536 => x"00000000",
    30537 => x"00000000", 30538 => x"00000000", 30539 => x"00000000",
    30540 => x"00000000", 30541 => x"00000000", 30542 => x"00000000",
    30543 => x"00000000", 30544 => x"00000000", 30545 => x"00000000",
    30546 => x"00000000", 30547 => x"00000000", 30548 => x"00000000",
    30549 => x"00000000", 30550 => x"00000000", 30551 => x"00000000",
    30552 => x"00000000", 30553 => x"00000000", 30554 => x"00000000",
    30555 => x"00000000", 30556 => x"00000000", 30557 => x"00000000",
    30558 => x"00000000", 30559 => x"00000000", 30560 => x"00000000",
    30561 => x"00000000", 30562 => x"00000000", 30563 => x"00000000",
    30564 => x"00000000", 30565 => x"00000000", 30566 => x"00000000",
    30567 => x"00000000", 30568 => x"00000000", 30569 => x"00000000",
    30570 => x"00000000", 30571 => x"00000000", 30572 => x"00000000",
    30573 => x"00000000", 30574 => x"00000000", 30575 => x"00000000",
    30576 => x"00000000", 30577 => x"00000000", 30578 => x"00000000",
    30579 => x"00000000", 30580 => x"00000000", 30581 => x"00000000",
    30582 => x"00000000", 30583 => x"00000000", 30584 => x"00000000",
    30585 => x"00000000", 30586 => x"00000000", 30587 => x"00000000",
    30588 => x"00000000", 30589 => x"00000000", 30590 => x"00000000",
    30591 => x"00000000", 30592 => x"00000000", 30593 => x"00000000",
    30594 => x"00000000", 30595 => x"00000000", 30596 => x"00000000",
    30597 => x"00000000", 30598 => x"00000000", 30599 => x"00000000",
    30600 => x"00000000", 30601 => x"00000000", 30602 => x"00000000",
    30603 => x"00000000", 30604 => x"00000000", 30605 => x"00000000",
    30606 => x"00000000", 30607 => x"00000000", 30608 => x"00000000",
    30609 => x"00000000", 30610 => x"00000000", 30611 => x"00000000",
    30612 => x"00000000", 30613 => x"00000000", 30614 => x"00000000",
    30615 => x"00000000", 30616 => x"00000000", 30617 => x"00000000",
    30618 => x"00000000", 30619 => x"00000000", 30620 => x"00000000",
    30621 => x"00000000", 30622 => x"00000000", 30623 => x"00000000",
    30624 => x"00000000", 30625 => x"00000000", 30626 => x"00000000",
    30627 => x"00000000", 30628 => x"00000000", 30629 => x"00000000",
    30630 => x"00000000", 30631 => x"00000000", 30632 => x"00000000",
    30633 => x"00000000", 30634 => x"00000000", 30635 => x"00000000",
    30636 => x"00000000", 30637 => x"00000000", 30638 => x"00000000",
    30639 => x"00000000", 30640 => x"00000000", 30641 => x"00000000",
    30642 => x"00000000", 30643 => x"00000000", 30644 => x"00000000",
    30645 => x"00000000", 30646 => x"00000000", 30647 => x"00000000",
    30648 => x"00000000", 30649 => x"00000000", 30650 => x"00000000",
    30651 => x"00000000", 30652 => x"00000000", 30653 => x"00000000",
    30654 => x"00000000", 30655 => x"00000000", 30656 => x"00000000",
    30657 => x"00000000", 30658 => x"00000000", 30659 => x"00000000",
    30660 => x"00000000", 30661 => x"00000000", 30662 => x"00000000",
    30663 => x"00000000", 30664 => x"00000000", 30665 => x"00000000",
    30666 => x"00000000", 30667 => x"00000000", 30668 => x"00000000",
    30669 => x"00000000", 30670 => x"00000000", 30671 => x"00000000",
    30672 => x"00000000", 30673 => x"00000000", 30674 => x"00000000",
    30675 => x"00000000", 30676 => x"00000000", 30677 => x"00000000",
    30678 => x"00000000", 30679 => x"00000000", 30680 => x"00000000",
    30681 => x"00000000", 30682 => x"00000000", 30683 => x"00000000",
    30684 => x"00000000", 30685 => x"00000000", 30686 => x"00000000",
    30687 => x"00000000", 30688 => x"00000000", 30689 => x"00000000",
    30690 => x"00000000", 30691 => x"00000000", 30692 => x"00000000",
    30693 => x"00000000", 30694 => x"00000000", 30695 => x"00000000",
    30696 => x"00000000", 30697 => x"00000000", 30698 => x"00000000",
    30699 => x"00000000", 30700 => x"00000000", 30701 => x"00000000",
    30702 => x"00000000", 30703 => x"00000000", 30704 => x"00000000",
    30705 => x"00000000", 30706 => x"00000000", 30707 => x"00000000",
    30708 => x"00000000", 30709 => x"00000000", 30710 => x"00000000",
    30711 => x"00000000", 30712 => x"00000000", 30713 => x"00000000",
    30714 => x"00000000", 30715 => x"00000000", 30716 => x"00000000",
    30717 => x"00000000", 30718 => x"00000000", 30719 => x"00000000",
    30720 => x"00000000", 30721 => x"00000000", 30722 => x"00000000",
    30723 => x"00000000", 30724 => x"00000000", 30725 => x"00000000",
    30726 => x"00000000", 30727 => x"00000000", 30728 => x"00000000",
    30729 => x"00000000", 30730 => x"00000000", 30731 => x"00000000",
    30732 => x"00000000", 30733 => x"00000000", 30734 => x"00000000",
    30735 => x"00000000", 30736 => x"00000000", 30737 => x"00000000",
    30738 => x"00000000", 30739 => x"00000000", 30740 => x"00000000",
    30741 => x"00000000", 30742 => x"00000000", 30743 => x"00000000",
    30744 => x"00000000", 30745 => x"00000000", 30746 => x"00000000",
    30747 => x"00000000", 30748 => x"00000000", 30749 => x"00000000",
    30750 => x"00000000", 30751 => x"00000000", 30752 => x"00000000",
    30753 => x"00000000", 30754 => x"00000000", 30755 => x"00000000",
    30756 => x"00000000", 30757 => x"00000000", 30758 => x"00000000",
    30759 => x"00000000", 30760 => x"00000000", 30761 => x"00000000",
    30762 => x"00000000", 30763 => x"00000000", 30764 => x"00000000",
    30765 => x"00000000", 30766 => x"00000000", 30767 => x"00000000",
    30768 => x"00000000", 30769 => x"00000000", 30770 => x"00000000",
    30771 => x"00000000", 30772 => x"00000000", 30773 => x"00000000",
    30774 => x"00000000", 30775 => x"00000000", 30776 => x"00000000",
    30777 => x"00000000", 30778 => x"00000000", 30779 => x"00000000",
    30780 => x"00000000", 30781 => x"00000000", 30782 => x"00000000",
    30783 => x"00000000", 30784 => x"00000000", 30785 => x"00000000",
    30786 => x"00000000", 30787 => x"00000000", 30788 => x"00000000",
    30789 => x"00000000", 30790 => x"00000000", 30791 => x"00000000",
    30792 => x"00000000", 30793 => x"00000000", 30794 => x"00000000",
    30795 => x"00000000", 30796 => x"00000000", 30797 => x"00000000",
    30798 => x"00000000", 30799 => x"00000000", 30800 => x"00000000",
    30801 => x"00000000", 30802 => x"00000000", 30803 => x"00000000",
    30804 => x"00000000", 30805 => x"00000000", 30806 => x"00000000",
    30807 => x"00000000", 30808 => x"00000000", 30809 => x"00000000",
    30810 => x"00000000", 30811 => x"00000000", 30812 => x"00000000",
    30813 => x"00000000", 30814 => x"00000000", 30815 => x"00000000",
    30816 => x"00000000", 30817 => x"00000000", 30818 => x"00000000",
    30819 => x"00000000", 30820 => x"00000000", 30821 => x"00000000",
    30822 => x"00000000", 30823 => x"00000000", 30824 => x"00000000",
    30825 => x"00000000", 30826 => x"00000000", 30827 => x"00000000",
    30828 => x"00000000", 30829 => x"00000000", 30830 => x"00000000",
    30831 => x"00000000", 30832 => x"00000000", 30833 => x"00000000",
    30834 => x"00000000", 30835 => x"00000000", 30836 => x"00000000",
    30837 => x"00000000", 30838 => x"00000000", 30839 => x"00000000",
    30840 => x"00000000", 30841 => x"00000000", 30842 => x"00000000",
    30843 => x"00000000", 30844 => x"00000000", 30845 => x"00000000",
    30846 => x"00000000", 30847 => x"00000000", 30848 => x"00000000",
    30849 => x"00000000", 30850 => x"00000000", 30851 => x"00000000",
    30852 => x"00000000", 30853 => x"00000000", 30854 => x"00000000",
    30855 => x"00000000", 30856 => x"00000000", 30857 => x"00000000",
    30858 => x"00000000", 30859 => x"00000000", 30860 => x"00000000",
    30861 => x"00000000", 30862 => x"00000000", 30863 => x"00000000",
    30864 => x"00000000", 30865 => x"00000000", 30866 => x"00000000",
    30867 => x"00000000", 30868 => x"00000000", 30869 => x"00000000",
    30870 => x"00000000", 30871 => x"00000000", 30872 => x"00000000",
    30873 => x"00000000", 30874 => x"00000000", 30875 => x"00000000",
    30876 => x"00000000", 30877 => x"00000000", 30878 => x"00000000",
    30879 => x"00000000", 30880 => x"00000000", 30881 => x"00000000",
    30882 => x"00000000", 30883 => x"00000000", 30884 => x"00000000",
    30885 => x"00000000", 30886 => x"00000000", 30887 => x"00000000",
    30888 => x"00000000", 30889 => x"00000000", 30890 => x"00000000",
    30891 => x"00000000", 30892 => x"00000000", 30893 => x"00000000",
    30894 => x"00000000", 30895 => x"00000000", 30896 => x"00000000",
    30897 => x"00000000", 30898 => x"00000000", 30899 => x"00000000",
    30900 => x"00000000", 30901 => x"00000000", 30902 => x"00000000",
    30903 => x"00000000", 30904 => x"00000000", 30905 => x"00000000",
    30906 => x"00000000", 30907 => x"00000000", 30908 => x"00000000",
    30909 => x"00000000", 30910 => x"00000000", 30911 => x"00000000",
    30912 => x"00000000", 30913 => x"00000000", 30914 => x"00000000",
    30915 => x"00000000", 30916 => x"00000000", 30917 => x"00000000",
    30918 => x"00000000", 30919 => x"00000000", 30920 => x"00000000",
    30921 => x"00000000", 30922 => x"00000000", 30923 => x"00000000",
    30924 => x"00000000", 30925 => x"00000000", 30926 => x"00000000",
    30927 => x"00000000", 30928 => x"00000000", 30929 => x"00000000",
    30930 => x"00000000", 30931 => x"00000000", 30932 => x"00000000",
    30933 => x"00000000", 30934 => x"00000000", 30935 => x"00000000",
    30936 => x"00000000", 30937 => x"00000000", 30938 => x"00000000",
    30939 => x"00000000", 30940 => x"00000000", 30941 => x"00000000",
    30942 => x"00000000", 30943 => x"00000000", 30944 => x"00000000",
    30945 => x"00000000", 30946 => x"00000000", 30947 => x"00000000",
    30948 => x"00000000", 30949 => x"00000000", 30950 => x"00000000",
    30951 => x"00000000", 30952 => x"00000000", 30953 => x"00000000",
    30954 => x"00000000", 30955 => x"00000000", 30956 => x"00000000",
    30957 => x"00000000", 30958 => x"00000000", 30959 => x"00000000",
    30960 => x"00000000", 30961 => x"00000000", 30962 => x"00000000",
    30963 => x"00000000", 30964 => x"00000000", 30965 => x"00000000",
    30966 => x"00000000", 30967 => x"00000000", 30968 => x"00000000",
    30969 => x"00000000", 30970 => x"00000000", 30971 => x"00000000",
    30972 => x"00000000", 30973 => x"00000000", 30974 => x"00000000",
    30975 => x"00000000", 30976 => x"00000000", 30977 => x"00000000",
    30978 => x"00000000", 30979 => x"00000000", 30980 => x"00000000",
    30981 => x"00000000", 30982 => x"00000000", 30983 => x"00000000",
    30984 => x"00000000", 30985 => x"00000000", 30986 => x"00000000",
    30987 => x"00000000", 30988 => x"00000000", 30989 => x"00000000",
    30990 => x"00000000", 30991 => x"00000000", 30992 => x"00000000",
    30993 => x"00000000", 30994 => x"00000000", 30995 => x"00000000",
    30996 => x"00000000", 30997 => x"00000000", 30998 => x"00000000",
    30999 => x"00000000", 31000 => x"00000000", 31001 => x"00000000",
    31002 => x"00000000", 31003 => x"00000000", 31004 => x"00000000",
    31005 => x"00000000", 31006 => x"00000000", 31007 => x"00000000",
    31008 => x"00000000", 31009 => x"00000000", 31010 => x"00000000",
    31011 => x"00000000", 31012 => x"00000000", 31013 => x"00000000",
    31014 => x"00000000", 31015 => x"00000000", 31016 => x"00000000",
    31017 => x"00000000", 31018 => x"00000000", 31019 => x"00000000",
    31020 => x"00000000", 31021 => x"00000000", 31022 => x"00000000",
    31023 => x"00000000", 31024 => x"00000000", 31025 => x"00000000",
    31026 => x"00000000", 31027 => x"00000000", 31028 => x"00000000",
    31029 => x"00000000", 31030 => x"00000000", 31031 => x"00000000",
    31032 => x"00000000", 31033 => x"00000000", 31034 => x"00000000",
    31035 => x"00000000", 31036 => x"00000000", 31037 => x"00000000",
    31038 => x"00000000", 31039 => x"00000000", 31040 => x"00000000",
    31041 => x"00000000", 31042 => x"00000000", 31043 => x"00000000",
    31044 => x"00000000", 31045 => x"00000000", 31046 => x"00000000",
    31047 => x"00000000", 31048 => x"00000000", 31049 => x"00000000",
    31050 => x"00000000", 31051 => x"00000000", 31052 => x"00000000",
    31053 => x"00000000", 31054 => x"00000000", 31055 => x"00000000",
    31056 => x"00000000", 31057 => x"00000000", 31058 => x"00000000",
    31059 => x"00000000", 31060 => x"00000000", 31061 => x"00000000",
    31062 => x"00000000", 31063 => x"00000000", 31064 => x"00000000",
    31065 => x"00000000", 31066 => x"00000000", 31067 => x"00000000",
    31068 => x"00000000", 31069 => x"00000000", 31070 => x"00000000",
    31071 => x"00000000", 31072 => x"00000000", 31073 => x"00000000",
    31074 => x"00000000", 31075 => x"00000000", 31076 => x"00000000",
    31077 => x"00000000", 31078 => x"00000000", 31079 => x"00000000",
    31080 => x"00000000", 31081 => x"00000000", 31082 => x"00000000",
    31083 => x"00000000", 31084 => x"00000000", 31085 => x"00000000",
    31086 => x"00000000", 31087 => x"00000000", 31088 => x"00000000",
    31089 => x"00000000", 31090 => x"00000000", 31091 => x"00000000",
    31092 => x"00000000", 31093 => x"00000000", 31094 => x"00000000",
    31095 => x"00000000", 31096 => x"00000000", 31097 => x"00000000",
    31098 => x"00000000", 31099 => x"00000000", 31100 => x"00000000",
    31101 => x"00000000", 31102 => x"00000000", 31103 => x"00000000",
    31104 => x"00000000", 31105 => x"00000000", 31106 => x"00000000",
    31107 => x"00000000", 31108 => x"00000000", 31109 => x"00000000",
    31110 => x"00000000", 31111 => x"00000000", 31112 => x"00000000",
    31113 => x"00000000", 31114 => x"00000000", 31115 => x"00000000",
    31116 => x"00000000", 31117 => x"00000000", 31118 => x"00000000",
    31119 => x"00000000", 31120 => x"00000000", 31121 => x"00000000",
    31122 => x"00000000", 31123 => x"00000000", 31124 => x"00000000",
    31125 => x"00000000", 31126 => x"00000000", 31127 => x"00000000",
    31128 => x"00000000", 31129 => x"00000000", 31130 => x"00000000",
    31131 => x"00000000", 31132 => x"00000000", 31133 => x"00000000",
    31134 => x"00000000", 31135 => x"00000000", 31136 => x"00000000",
    31137 => x"00000000", 31138 => x"00000000", 31139 => x"00000000",
    31140 => x"00000000", 31141 => x"00000000", 31142 => x"00000000",
    31143 => x"00000000", 31144 => x"00000000", 31145 => x"00000000",
    31146 => x"00000000", 31147 => x"00000000", 31148 => x"00000000",
    31149 => x"00000000", 31150 => x"00000000", 31151 => x"00000000",
    31152 => x"00000000", 31153 => x"00000000", 31154 => x"00000000",
    31155 => x"00000000", 31156 => x"00000000", 31157 => x"00000000",
    31158 => x"00000000", 31159 => x"00000000", 31160 => x"00000000",
    31161 => x"00000000", 31162 => x"00000000", 31163 => x"00000000",
    31164 => x"00000000", 31165 => x"00000000", 31166 => x"00000000",
    31167 => x"00000000", 31168 => x"00000000", 31169 => x"00000000",
    31170 => x"00000000", 31171 => x"00000000", 31172 => x"00000000",
    31173 => x"00000000", 31174 => x"00000000", 31175 => x"00000000",
    31176 => x"00000000", 31177 => x"00000000", 31178 => x"00000000",
    31179 => x"00000000", 31180 => x"00000000", 31181 => x"00000000",
    31182 => x"00000000", 31183 => x"00000000", 31184 => x"00000000",
    31185 => x"00000000", 31186 => x"00000000", 31187 => x"00000000",
    31188 => x"00000000", 31189 => x"00000000", 31190 => x"00000000",
    31191 => x"00000000", 31192 => x"00000000", 31193 => x"00000000",
    31194 => x"00000000", 31195 => x"00000000", 31196 => x"00000000",
    31197 => x"00000000", 31198 => x"00000000", 31199 => x"00000000",
    31200 => x"00000000", 31201 => x"00000000", 31202 => x"00000000",
    31203 => x"00000000", 31204 => x"00000000", 31205 => x"00000000",
    31206 => x"00000000", 31207 => x"00000000", 31208 => x"00000000",
    31209 => x"00000000", 31210 => x"00000000", 31211 => x"00000000",
    31212 => x"00000000", 31213 => x"00000000", 31214 => x"00000000",
    31215 => x"00000000", 31216 => x"00000000", 31217 => x"00000000",
    31218 => x"00000000", 31219 => x"00000000", 31220 => x"00000000",
    31221 => x"00000000", 31222 => x"00000000", 31223 => x"00000000",
    31224 => x"00000000", 31225 => x"00000000", 31226 => x"00000000",
    31227 => x"00000000", 31228 => x"00000000", 31229 => x"00000000",
    31230 => x"00000000", 31231 => x"00000000", 31232 => x"00000000",
    31233 => x"00000000", 31234 => x"00000000", 31235 => x"00000000",
    31236 => x"00000000", 31237 => x"00000000", 31238 => x"00000000",
    31239 => x"00000000", 31240 => x"00000000", 31241 => x"00000000",
    31242 => x"00000000", 31243 => x"00000000", 31244 => x"00000000",
    31245 => x"00000000", 31246 => x"00000000", 31247 => x"00000000",
    31248 => x"00000000", 31249 => x"00000000", 31250 => x"00000000",
    31251 => x"00000000", 31252 => x"00000000", 31253 => x"00000000",
    31254 => x"00000000", 31255 => x"00000000", 31256 => x"00000000",
    31257 => x"00000000", 31258 => x"00000000", 31259 => x"00000000",
    31260 => x"00000000", 31261 => x"00000000", 31262 => x"00000000",
    31263 => x"00000000", 31264 => x"00000000", 31265 => x"00000000",
    31266 => x"00000000", 31267 => x"00000000", 31268 => x"00000000",
    31269 => x"00000000", 31270 => x"00000000", 31271 => x"00000000",
    31272 => x"00000000", 31273 => x"00000000", 31274 => x"00000000",
    31275 => x"00000000", 31276 => x"00000000", 31277 => x"00000000",
    31278 => x"00000000", 31279 => x"00000000", 31280 => x"00000000",
    31281 => x"00000000", 31282 => x"00000000", 31283 => x"00000000",
    31284 => x"00000000", 31285 => x"00000000", 31286 => x"00000000",
    31287 => x"00000000", 31288 => x"00000000", 31289 => x"00000000",
    31290 => x"00000000", 31291 => x"00000000", 31292 => x"00000000",
    31293 => x"00000000", 31294 => x"00000000", 31295 => x"00000000",
    31296 => x"00000000", 31297 => x"00000000", 31298 => x"00000000",
    31299 => x"00000000", 31300 => x"00000000", 31301 => x"00000000",
    31302 => x"00000000", 31303 => x"00000000", 31304 => x"00000000",
    31305 => x"00000000", 31306 => x"00000000", 31307 => x"00000000",
    31308 => x"00000000", 31309 => x"00000000", 31310 => x"00000000",
    31311 => x"00000000", 31312 => x"00000000", 31313 => x"00000000",
    31314 => x"00000000", 31315 => x"00000000", 31316 => x"00000000",
    31317 => x"00000000", 31318 => x"00000000", 31319 => x"00000000",
    31320 => x"00000000", 31321 => x"00000000", 31322 => x"00000000",
    31323 => x"00000000", 31324 => x"00000000", 31325 => x"00000000",
    31326 => x"00000000", 31327 => x"00000000", 31328 => x"00000000",
    31329 => x"00000000", 31330 => x"00000000", 31331 => x"00000000",
    31332 => x"00000000", 31333 => x"00000000", 31334 => x"00000000",
    31335 => x"00000000", 31336 => x"00000000", 31337 => x"00000000",
    31338 => x"00000000", 31339 => x"00000000", 31340 => x"00000000",
    31341 => x"00000000", 31342 => x"00000000", 31343 => x"00000000",
    31344 => x"00000000", 31345 => x"00000000", 31346 => x"00000000",
    31347 => x"00000000", 31348 => x"00000000", 31349 => x"00000000",
    31350 => x"00000000", 31351 => x"00000000", 31352 => x"00000000",
    31353 => x"00000000", 31354 => x"00000000", 31355 => x"00000000",
    31356 => x"00000000", 31357 => x"00000000", 31358 => x"00000000",
    31359 => x"00000000", 31360 => x"00000000", 31361 => x"00000000",
    31362 => x"00000000", 31363 => x"00000000", 31364 => x"00000000",
    31365 => x"00000000", 31366 => x"00000000", 31367 => x"00000000",
    31368 => x"00000000", 31369 => x"00000000", 31370 => x"00000000",
    31371 => x"00000000", 31372 => x"00000000", 31373 => x"00000000",
    31374 => x"00000000", 31375 => x"00000000", 31376 => x"00000000",
    31377 => x"00000000", 31378 => x"00000000", 31379 => x"00000000",
    31380 => x"00000000", 31381 => x"00000000", 31382 => x"00000000",
    31383 => x"00000000", 31384 => x"00000000", 31385 => x"00000000",
    31386 => x"00000000", 31387 => x"00000000", 31388 => x"00000000",
    31389 => x"00000000", 31390 => x"00000000", 31391 => x"00000000",
    31392 => x"00000000", 31393 => x"00000000", 31394 => x"00000000",
    31395 => x"00000000", 31396 => x"00000000", 31397 => x"00000000",
    31398 => x"00000000", 31399 => x"00000000", 31400 => x"00000000",
    31401 => x"00000000", 31402 => x"00000000", 31403 => x"00000000",
    31404 => x"00000000", 31405 => x"00000000", 31406 => x"00000000",
    31407 => x"00000000", 31408 => x"00000000", 31409 => x"00000000",
    31410 => x"00000000", 31411 => x"00000000", 31412 => x"00000000",
    31413 => x"00000000", 31414 => x"00000000", 31415 => x"00000000",
    31416 => x"00000000", 31417 => x"00000000", 31418 => x"00000000",
    31419 => x"00000000", 31420 => x"00000000", 31421 => x"00000000",
    31422 => x"00000000", 31423 => x"00000000", 31424 => x"00000000",
    31425 => x"00000000", 31426 => x"00000000", 31427 => x"00000000",
    31428 => x"00000000", 31429 => x"00000000", 31430 => x"00000000",
    31431 => x"00000000", 31432 => x"00000000", 31433 => x"00000000",
    31434 => x"00000000", 31435 => x"00000000", 31436 => x"00000000",
    31437 => x"00000000", 31438 => x"00000000", 31439 => x"00000000",
    31440 => x"00000000", 31441 => x"00000000", 31442 => x"00000000",
    31443 => x"00000000", 31444 => x"00000000", 31445 => x"00000000",
    31446 => x"00000000", 31447 => x"00000000", 31448 => x"00000000",
    31449 => x"00000000", 31450 => x"00000000", 31451 => x"00000000",
    31452 => x"00000000", 31453 => x"00000000", 31454 => x"00000000",
    31455 => x"00000000", 31456 => x"00000000", 31457 => x"00000000",
    31458 => x"00000000", 31459 => x"00000000", 31460 => x"00000000",
    31461 => x"00000000", 31462 => x"00000000", 31463 => x"00000000",
    31464 => x"00000000", 31465 => x"00000000", 31466 => x"00000000",
    31467 => x"00000000", 31468 => x"00000000", 31469 => x"00000000",
    31470 => x"00000000", 31471 => x"00000000", 31472 => x"00000000",
    31473 => x"00000000", 31474 => x"00000000", 31475 => x"00000000",
    31476 => x"00000000", 31477 => x"00000000", 31478 => x"00000000",
    31479 => x"00000000", 31480 => x"00000000", 31481 => x"00000000",
    31482 => x"00000000", 31483 => x"00000000", 31484 => x"00000000",
    31485 => x"00000000", 31486 => x"00000000", 31487 => x"00000000",
    31488 => x"00000000", 31489 => x"00000000", 31490 => x"00000000",
    31491 => x"00000000", 31492 => x"00000000", 31493 => x"00000000",
    31494 => x"00000000", 31495 => x"00000000", 31496 => x"00000000",
    31497 => x"00000000", 31498 => x"00000000", 31499 => x"00000000",
    31500 => x"00000000", 31501 => x"00000000", 31502 => x"00000000",
    31503 => x"00000000", 31504 => x"00000000", 31505 => x"00000000",
    31506 => x"00000000", 31507 => x"00000000", 31508 => x"00000000",
    31509 => x"00000000", 31510 => x"00000000", 31511 => x"00000000",
    31512 => x"00000000", 31513 => x"00000000", 31514 => x"00000000",
    31515 => x"00000000", 31516 => x"00000000", 31517 => x"00000000",
    31518 => x"00000000", 31519 => x"00000000", 31520 => x"00000000",
    31521 => x"00000000", 31522 => x"00000000", 31523 => x"00000000",
    31524 => x"00000000", 31525 => x"00000000", 31526 => x"00000000",
    31527 => x"00000000", 31528 => x"00000000", 31529 => x"00000000",
    31530 => x"00000000", 31531 => x"00000000", 31532 => x"00000000",
    31533 => x"00000000", 31534 => x"00000000", 31535 => x"00000000",
    31536 => x"00000000", 31537 => x"00000000", 31538 => x"00000000",
    31539 => x"00000000", 31540 => x"00000000", 31541 => x"00000000",
    31542 => x"00000000", 31543 => x"00000000", 31544 => x"00000000",
    31545 => x"00000000", 31546 => x"00000000", 31547 => x"00000000",
    31548 => x"00000000", 31549 => x"00000000", 31550 => x"00000000",
    31551 => x"00000000", 31552 => x"00000000", 31553 => x"00000000",
    31554 => x"00000000", 31555 => x"00000000", 31556 => x"00000000",
    31557 => x"00000000", 31558 => x"00000000", 31559 => x"00000000",
    31560 => x"00000000", 31561 => x"00000000", 31562 => x"00000000",
    31563 => x"00000000", 31564 => x"00000000", 31565 => x"00000000",
    31566 => x"00000000", 31567 => x"00000000", 31568 => x"00000000",
    31569 => x"00000000", 31570 => x"00000000", 31571 => x"00000000",
    31572 => x"00000000", 31573 => x"00000000", 31574 => x"00000000",
    31575 => x"00000000", 31576 => x"00000000", 31577 => x"00000000",
    31578 => x"00000000", 31579 => x"00000000", 31580 => x"00000000",
    31581 => x"00000000", 31582 => x"00000000", 31583 => x"00000000",
    31584 => x"00000000", 31585 => x"00000000", 31586 => x"00000000",
    31587 => x"00000000", 31588 => x"00000000", 31589 => x"00000000",
    31590 => x"00000000", 31591 => x"00000000", 31592 => x"00000000",
    31593 => x"00000000", 31594 => x"00000000", 31595 => x"00000000",
    31596 => x"00000000", 31597 => x"00000000", 31598 => x"00000000",
    31599 => x"00000000", 31600 => x"00000000", 31601 => x"00000000",
    31602 => x"00000000", 31603 => x"00000000", 31604 => x"00000000",
    31605 => x"00000000", 31606 => x"00000000", 31607 => x"00000000",
    31608 => x"00000000", 31609 => x"00000000", 31610 => x"00000000",
    31611 => x"00000000", 31612 => x"00000000", 31613 => x"00000000",
    31614 => x"00000000", 31615 => x"00000000", 31616 => x"00000000",
    31617 => x"00000000", 31618 => x"00000000", 31619 => x"00000000",
    31620 => x"00000000", 31621 => x"00000000", 31622 => x"00000000",
    31623 => x"00000000", 31624 => x"00000000", 31625 => x"00000000",
    31626 => x"00000000", 31627 => x"00000000", 31628 => x"00000000",
    31629 => x"00000000", 31630 => x"00000000", 31631 => x"00000000",
    31632 => x"00000000", 31633 => x"00000000", 31634 => x"00000000",
    31635 => x"00000000", 31636 => x"00000000", 31637 => x"00000000",
    31638 => x"00000000", 31639 => x"00000000", 31640 => x"00000000",
    31641 => x"00000000", 31642 => x"00000000", 31643 => x"00000000",
    31644 => x"00000000", 31645 => x"00000000", 31646 => x"00000000",
    31647 => x"00000000", 31648 => x"00000000", 31649 => x"00000000",
    31650 => x"00000000", 31651 => x"00000000", 31652 => x"00000000",
    31653 => x"00000000", 31654 => x"00000000", 31655 => x"00000000",
    31656 => x"00000000", 31657 => x"00000000", 31658 => x"00000000",
    31659 => x"00000000", 31660 => x"00000000", 31661 => x"00000000",
    31662 => x"00000000", 31663 => x"00000000", 31664 => x"00000000",
    31665 => x"00000000", 31666 => x"00000000", 31667 => x"00000000",
    31668 => x"00000000", 31669 => x"00000000", 31670 => x"00000000",
    31671 => x"00000000", 31672 => x"00000000", 31673 => x"00000000",
    31674 => x"00000000", 31675 => x"00000000", 31676 => x"00000000",
    31677 => x"00000000", 31678 => x"00000000", 31679 => x"00000000",
    31680 => x"00000000", 31681 => x"00000000", 31682 => x"00000000",
    31683 => x"00000000", 31684 => x"00000000", 31685 => x"00000000",
    31686 => x"00000000", 31687 => x"00000000", 31688 => x"00000000",
    31689 => x"00000000", 31690 => x"00000000", 31691 => x"00000000",
    31692 => x"00000000", 31693 => x"00000000", 31694 => x"00000000",
    31695 => x"00000000", 31696 => x"00000000", 31697 => x"00000000",
    31698 => x"00000000", 31699 => x"00000000", 31700 => x"00000000",
    31701 => x"00000000", 31702 => x"00000000", 31703 => x"00000000",
    31704 => x"00000000", 31705 => x"00000000", 31706 => x"00000000",
    31707 => x"00000000", 31708 => x"00000000", 31709 => x"00000000",
    31710 => x"00000000", 31711 => x"00000000", 31712 => x"00000000",
    31713 => x"00000000", 31714 => x"00000000", 31715 => x"00000000",
    31716 => x"00000000", 31717 => x"00000000", 31718 => x"00000000",
    31719 => x"00000000", 31720 => x"00000000", 31721 => x"00000000",
    31722 => x"00000000", 31723 => x"00000000", 31724 => x"00000000",
    31725 => x"00000000", 31726 => x"00000000", 31727 => x"00000000",
    31728 => x"00000000", 31729 => x"00000000", 31730 => x"00000000",
    31731 => x"00000000", 31732 => x"00000000", 31733 => x"00000000",
    31734 => x"00000000", 31735 => x"00000000", 31736 => x"00000000",
    31737 => x"00000000", 31738 => x"00000000", 31739 => x"00000000",
    31740 => x"00000000", 31741 => x"00000000", 31742 => x"00000000",
    31743 => x"00000000", 31744 => x"00000000", 31745 => x"00000000",
    31746 => x"00000000", 31747 => x"00000000", 31748 => x"00000000",
    31749 => x"00000000", 31750 => x"00000000", 31751 => x"00000000",
    31752 => x"00000000", 31753 => x"00000000", 31754 => x"00000000",
    31755 => x"00000000", 31756 => x"00000000", 31757 => x"00000000",
    31758 => x"00000000", 31759 => x"00000000", 31760 => x"00000000",
    31761 => x"00000000", 31762 => x"00000000", 31763 => x"00000000",
    31764 => x"00000000", 31765 => x"00000000", 31766 => x"00000000",
    31767 => x"00000000", 31768 => x"00000000", 31769 => x"00000000",
    31770 => x"00000000", 31771 => x"00000000", 31772 => x"00000000",
    31773 => x"00000000", 31774 => x"00000000", 31775 => x"00000000",
    31776 => x"00000000", 31777 => x"00000000", 31778 => x"00000000",
    31779 => x"00000000", 31780 => x"00000000", 31781 => x"00000000",
    31782 => x"00000000", 31783 => x"00000000", 31784 => x"00000000",
    31785 => x"00000000", 31786 => x"00000000", 31787 => x"00000000",
    31788 => x"00000000", 31789 => x"00000000", 31790 => x"00000000",
    31791 => x"00000000", 31792 => x"00000000", 31793 => x"00000000",
    31794 => x"00000000", 31795 => x"00000000", 31796 => x"00000000",
    31797 => x"00000000", 31798 => x"00000000", 31799 => x"00000000",
    31800 => x"00000000", 31801 => x"00000000", 31802 => x"00000000",
    31803 => x"00000000", 31804 => x"00000000", 31805 => x"00000000",
    31806 => x"00000000", 31807 => x"00000000", 31808 => x"00000000",
    31809 => x"00000000", 31810 => x"00000000", 31811 => x"00000000",
    31812 => x"00000000", 31813 => x"00000000", 31814 => x"00000000",
    31815 => x"00000000", 31816 => x"00000000", 31817 => x"00000000",
    31818 => x"00000000", 31819 => x"00000000", 31820 => x"00000000",
    31821 => x"00000000", 31822 => x"00000000", 31823 => x"00000000",
    31824 => x"00000000", 31825 => x"00000000", 31826 => x"00000000",
    31827 => x"00000000", 31828 => x"00000000", 31829 => x"00000000",
    31830 => x"00000000", 31831 => x"00000000", 31832 => x"00000000",
    31833 => x"00000000", 31834 => x"00000000", 31835 => x"00000000",
    31836 => x"00000000", 31837 => x"00000000", 31838 => x"00000000",
    31839 => x"00000000", 31840 => x"00000000", 31841 => x"00000000",
    31842 => x"00000000", 31843 => x"00000000", 31844 => x"00000000",
    31845 => x"00000000", 31846 => x"00000000", 31847 => x"00000000",
    31848 => x"00000000", 31849 => x"00000000", 31850 => x"00000000",
    31851 => x"00000000", 31852 => x"00000000", 31853 => x"00000000",
    31854 => x"00000000", 31855 => x"00000000", 31856 => x"00000000",
    31857 => x"00000000", 31858 => x"00000000", 31859 => x"00000000",
    31860 => x"00000000", 31861 => x"00000000", 31862 => x"00000000",
    31863 => x"00000000", 31864 => x"00000000", 31865 => x"00000000",
    31866 => x"00000000", 31867 => x"00000000", 31868 => x"00000000",
    31869 => x"00000000", 31870 => x"00000000", 31871 => x"00000000",
    31872 => x"00000000", 31873 => x"00000000", 31874 => x"00000000",
    31875 => x"00000000", 31876 => x"00000000", 31877 => x"00000000",
    31878 => x"00000000", 31879 => x"00000000", 31880 => x"00000000",
    31881 => x"00000000", 31882 => x"00000000", 31883 => x"00000000",
    31884 => x"00000000", 31885 => x"00000000", 31886 => x"00000000",
    31887 => x"00000000", 31888 => x"00000000", 31889 => x"00000000",
    31890 => x"00000000", 31891 => x"00000000", 31892 => x"00000000",
    31893 => x"00000000", 31894 => x"00000000", 31895 => x"00000000",
    31896 => x"00000000", 31897 => x"00000000", 31898 => x"00000000",
    31899 => x"00000000", 31900 => x"00000000", 31901 => x"00000000",
    31902 => x"00000000", 31903 => x"00000000", 31904 => x"00000000",
    31905 => x"00000000", 31906 => x"00000000", 31907 => x"00000000",
    31908 => x"00000000", 31909 => x"00000000", 31910 => x"00000000",
    31911 => x"00000000", 31912 => x"00000000", 31913 => x"00000000",
    31914 => x"00000000", 31915 => x"00000000", 31916 => x"00000000",
    31917 => x"00000000", 31918 => x"00000000", 31919 => x"00000000",
    31920 => x"00000000", 31921 => x"00000000", 31922 => x"00000000",
    31923 => x"00000000", 31924 => x"00000000", 31925 => x"00000000",
    31926 => x"00000000", 31927 => x"00000000", 31928 => x"00000000",
    31929 => x"00000000", 31930 => x"00000000", 31931 => x"00000000",
    31932 => x"00000000", 31933 => x"00000000", 31934 => x"00000000",
    31935 => x"00000000", 31936 => x"00000000", 31937 => x"00000000",
    31938 => x"00000000", 31939 => x"00000000", 31940 => x"00000000",
    31941 => x"00000000", 31942 => x"00000000", 31943 => x"00000000",
    31944 => x"00000000", 31945 => x"00000000", 31946 => x"00000000",
    31947 => x"00000000", 31948 => x"00000000", 31949 => x"00000000",
    31950 => x"00000000", 31951 => x"00000000", 31952 => x"00000000",
    31953 => x"00000000", 31954 => x"00000000", 31955 => x"00000000",
    31956 => x"00000000", 31957 => x"00000000", 31958 => x"00000000",
    31959 => x"00000000", 31960 => x"00000000", 31961 => x"00000000",
    31962 => x"00000000", 31963 => x"00000000", 31964 => x"00000000",
    31965 => x"00000000", 31966 => x"00000000", 31967 => x"00000000",
    31968 => x"00000000", 31969 => x"00000000", 31970 => x"00000000",
    31971 => x"00000000", 31972 => x"00000000", 31973 => x"00000000",
    31974 => x"00000000", 31975 => x"00000000", 31976 => x"00000000",
    31977 => x"00000000", 31978 => x"00000000", 31979 => x"00000000",
    31980 => x"00000000", 31981 => x"00000000", 31982 => x"00000000",
    31983 => x"00000000", 31984 => x"00000000", 31985 => x"00000000",
    31986 => x"00000000", 31987 => x"00000000", 31988 => x"00000000",
    31989 => x"00000000", 31990 => x"00000000", 31991 => x"00000000",
    31992 => x"00000000", 31993 => x"00000000", 31994 => x"00000000",
    31995 => x"00000000", 31996 => x"00000000", 31997 => x"00000000",
    31998 => x"00000000", 31999 => x"00000000", 32000 => x"00000000",
    32001 => x"00000000", 32002 => x"00000000", 32003 => x"00000000",
    32004 => x"00000000", 32005 => x"00000000", 32006 => x"00000000",
    32007 => x"00000000", 32008 => x"00000000", 32009 => x"00000000",
    32010 => x"00000000", 32011 => x"00000000", 32012 => x"00000000",
    32013 => x"00000000", 32014 => x"00000000", 32015 => x"00000000",
    32016 => x"00000000", 32017 => x"00000000", 32018 => x"00000000",
    32019 => x"00000000", 32020 => x"00000000", 32021 => x"00000000",
    32022 => x"00000000", 32023 => x"00000000", 32024 => x"00000000",
    32025 => x"00000000", 32026 => x"00000000", 32027 => x"00000000",
    32028 => x"00000000", 32029 => x"00000000", 32030 => x"00000000",
    32031 => x"00000000", 32032 => x"00000000", 32033 => x"00000000",
    32034 => x"00000000", 32035 => x"00000000", 32036 => x"00000000",
    32037 => x"00000000", 32038 => x"00000000", 32039 => x"00000000",
    32040 => x"00000000", 32041 => x"00000000", 32042 => x"00000000",
    32043 => x"00000000", 32044 => x"00000000", 32045 => x"00000000",
    32046 => x"00000000", 32047 => x"00000000", 32048 => x"00000000",
    32049 => x"00000000", 32050 => x"00000000", 32051 => x"00000000",
    32052 => x"00000000", 32053 => x"00000000", 32054 => x"00000000",
    32055 => x"00000000", 32056 => x"00000000", 32057 => x"00000000",
    32058 => x"00000000", 32059 => x"00000000", 32060 => x"00000000",
    32061 => x"00000000", 32062 => x"00000000", 32063 => x"00000000",
    32064 => x"00000000", 32065 => x"00000000", 32066 => x"00000000",
    32067 => x"00000000", 32068 => x"00000000", 32069 => x"00000000",
    32070 => x"00000000", 32071 => x"00000000", 32072 => x"00000000",
    32073 => x"00000000", 32074 => x"00000000", 32075 => x"00000000",
    32076 => x"00000000", 32077 => x"00000000", 32078 => x"00000000",
    32079 => x"00000000", 32080 => x"00000000", 32081 => x"00000000",
    32082 => x"00000000", 32083 => x"00000000", 32084 => x"00000000",
    32085 => x"00000000", 32086 => x"00000000", 32087 => x"00000000",
    32088 => x"00000000", 32089 => x"00000000", 32090 => x"00000000",
    32091 => x"00000000", 32092 => x"00000000", 32093 => x"00000000",
    32094 => x"00000000", 32095 => x"00000000", 32096 => x"00000000",
    32097 => x"00000000", 32098 => x"00000000", 32099 => x"00000000",
    32100 => x"00000000", 32101 => x"00000000", 32102 => x"00000000",
    32103 => x"00000000", 32104 => x"00000000", 32105 => x"00000000",
    32106 => x"00000000", 32107 => x"00000000", 32108 => x"00000000",
    32109 => x"00000000", 32110 => x"00000000", 32111 => x"00000000",
    32112 => x"00000000", 32113 => x"00000000", 32114 => x"00000000",
    32115 => x"00000000", 32116 => x"00000000", 32117 => x"00000000",
    32118 => x"00000000", 32119 => x"00000000", 32120 => x"00000000",
    32121 => x"00000000", 32122 => x"00000000", 32123 => x"00000000",
    32124 => x"00000000", 32125 => x"00000000", 32126 => x"00000000",
    32127 => x"00000000", 32128 => x"00000000", 32129 => x"00000000",
    32130 => x"00000000", 32131 => x"00000000", 32132 => x"00000000",
    32133 => x"00000000", 32134 => x"00000000", 32135 => x"00000000",
    32136 => x"00000000", 32137 => x"00000000", 32138 => x"00000000",
    32139 => x"00000000", 32140 => x"00000000", 32141 => x"00000000",
    32142 => x"00000000", 32143 => x"00000000", 32144 => x"00000000",
    32145 => x"00000000", 32146 => x"00000000", 32147 => x"00000000",
    32148 => x"00000000", 32149 => x"00000000", 32150 => x"00000000",
    32151 => x"00000000", 32152 => x"00000000", 32153 => x"00000000",
    32154 => x"00000000", 32155 => x"00000000", 32156 => x"00000000",
    32157 => x"00000000", 32158 => x"00000000", 32159 => x"00000000",
    32160 => x"00000000", 32161 => x"00000000", 32162 => x"00000000",
    32163 => x"00000000", 32164 => x"00000000", 32165 => x"00000000",
    32166 => x"00000000", 32167 => x"00000000", 32168 => x"00000000",
    32169 => x"00000000", 32170 => x"00000000", 32171 => x"00000000",
    32172 => x"00000000", 32173 => x"00000000", 32174 => x"00000000",
    32175 => x"00000000", 32176 => x"00000000", 32177 => x"00000000",
    32178 => x"00000000", 32179 => x"00000000", 32180 => x"00000000",
    32181 => x"00000000", 32182 => x"00000000", 32183 => x"00000000",
    32184 => x"00000000", 32185 => x"00000000", 32186 => x"00000000",
    32187 => x"00000000", 32188 => x"00000000", 32189 => x"00000000",
    32190 => x"00000000", 32191 => x"00000000", 32192 => x"00000000",
    32193 => x"00000000", 32194 => x"00000000", 32195 => x"00000000",
    32196 => x"00000000", 32197 => x"00000000", 32198 => x"00000000",
    32199 => x"00000000", 32200 => x"00000000", 32201 => x"00000000",
    32202 => x"00000000", 32203 => x"00000000", 32204 => x"00000000",
    32205 => x"00000000", 32206 => x"00000000", 32207 => x"00000000",
    32208 => x"00000000", 32209 => x"00000000", 32210 => x"00000000",
    32211 => x"00000000", 32212 => x"00000000", 32213 => x"00000000",
    32214 => x"00000000", 32215 => x"00000000", 32216 => x"00000000",
    32217 => x"00000000", 32218 => x"00000000", 32219 => x"00000000",
    32220 => x"00000000", 32221 => x"00000000", 32222 => x"00000000",
    32223 => x"00000000", 32224 => x"00000000", 32225 => x"00000000",
    32226 => x"00000000", 32227 => x"00000000", 32228 => x"00000000",
    32229 => x"00000000", 32230 => x"00000000", 32231 => x"00000000",
    32232 => x"00000000", 32233 => x"00000000", 32234 => x"00000000",
    32235 => x"00000000", 32236 => x"00000000", 32237 => x"00000000",
    32238 => x"00000000", 32239 => x"00000000", 32240 => x"00000000",
    32241 => x"00000000", 32242 => x"00000000", 32243 => x"00000000",
    32244 => x"00000000", 32245 => x"00000000", 32246 => x"00000000",
    32247 => x"00000000", 32248 => x"00000000", 32249 => x"00000000",
    32250 => x"00000000", 32251 => x"00000000", 32252 => x"00000000",
    32253 => x"00000000", 32254 => x"00000000", 32255 => x"00000000",
    32256 => x"00000000", 32257 => x"00000000", 32258 => x"00000000",
    32259 => x"00000000", 32260 => x"00000000", 32261 => x"00000000",
    32262 => x"00000000", 32263 => x"00000000", 32264 => x"00000000",
    32265 => x"00000000", 32266 => x"00000000", 32267 => x"00000000",
    32268 => x"00000000", 32269 => x"00000000", 32270 => x"00000000",
    32271 => x"00000000", 32272 => x"00000000", 32273 => x"00000000",
    32274 => x"00000000", 32275 => x"00000000", 32276 => x"00000000",
    32277 => x"00000000", 32278 => x"00000000", 32279 => x"00000000",
    32280 => x"00000000", 32281 => x"00000000", 32282 => x"00000000",
    32283 => x"00000000", 32284 => x"00000000", 32285 => x"00000000",
    32286 => x"00000000", 32287 => x"00000000", 32288 => x"00000000",
    32289 => x"00000000", 32290 => x"00000000", 32291 => x"00000000",
    32292 => x"00000000", 32293 => x"00000000", 32294 => x"00000000",
    32295 => x"00000000", 32296 => x"00000000", 32297 => x"00000000",
    32298 => x"00000000", 32299 => x"00000000", 32300 => x"00000000",
    32301 => x"00000000", 32302 => x"00000000", 32303 => x"00000000",
    32304 => x"00000000", 32305 => x"00000000", 32306 => x"00000000",
    32307 => x"00000000", 32308 => x"00000000", 32309 => x"00000000",
    32310 => x"00000000", 32311 => x"00000000", 32312 => x"00000000",
    32313 => x"00000000", 32314 => x"00000000", 32315 => x"00000000",
    32316 => x"00000000", 32317 => x"00000000", 32318 => x"00000000",
    32319 => x"00000000", 32320 => x"00000000", 32321 => x"00000000",
    32322 => x"00000000", 32323 => x"00000000", 32324 => x"00000000",
    32325 => x"00000000", 32326 => x"00000000", 32327 => x"00000000",
    32328 => x"00000000", 32329 => x"00000000", 32330 => x"00000000",
    32331 => x"00000000", 32332 => x"00000000", 32333 => x"00000000",
    32334 => x"00000000", 32335 => x"00000000", 32336 => x"00000000",
    32337 => x"00000000", 32338 => x"00000000", 32339 => x"00000000",
    32340 => x"00000000", 32341 => x"00000000", 32342 => x"00000000",
    32343 => x"00000000", 32344 => x"00000000", 32345 => x"00000000",
    32346 => x"00000000", 32347 => x"00000000", 32348 => x"00000000",
    32349 => x"00000000", 32350 => x"00000000", 32351 => x"00000000",
    32352 => x"00000000", 32353 => x"00000000", 32354 => x"00000000",
    32355 => x"00000000", 32356 => x"00000000", 32357 => x"00000000",
    32358 => x"00000000", 32359 => x"00000000", 32360 => x"00000000",
    32361 => x"00000000", 32362 => x"00000000", 32363 => x"00000000",
    32364 => x"00000000", 32365 => x"00000000", 32366 => x"00000000",
    32367 => x"00000000", 32368 => x"00000000", 32369 => x"00000000",
    32370 => x"00000000", 32371 => x"00000000", 32372 => x"00000000",
    32373 => x"00000000", 32374 => x"00000000", 32375 => x"00000000",
    32376 => x"00000000", 32377 => x"00000000", 32378 => x"00000000",
    32379 => x"00000000", 32380 => x"00000000", 32381 => x"00000000",
    32382 => x"00000000", 32383 => x"00000000", 32384 => x"00000000",
    32385 => x"00000000", 32386 => x"00000000", 32387 => x"00000000",
    32388 => x"00000000", 32389 => x"00000000", 32390 => x"00000000",
    32391 => x"00000000", 32392 => x"00000000", 32393 => x"00000000",
    32394 => x"00000000", 32395 => x"00000000", 32396 => x"00000000",
    32397 => x"00000000", 32398 => x"00000000", 32399 => x"00000000",
    32400 => x"00000000", 32401 => x"00000000", 32402 => x"00000000",
    32403 => x"00000000", 32404 => x"00000000", 32405 => x"00000000",
    32406 => x"00000000", 32407 => x"00000000", 32408 => x"00000000",
    32409 => x"00000000", 32410 => x"00000000", 32411 => x"00000000",
    32412 => x"00000000", 32413 => x"00000000", 32414 => x"00000000",
    32415 => x"00000000", 32416 => x"00000000", 32417 => x"00000000",
    32418 => x"00000000", 32419 => x"00000000", 32420 => x"00000000",
    32421 => x"00000000", 32422 => x"00000000", 32423 => x"00000000",
    32424 => x"00000000", 32425 => x"00000000", 32426 => x"00000000",
    32427 => x"00000000", 32428 => x"00000000", 32429 => x"00000000",
    32430 => x"00000000", 32431 => x"00000000", 32432 => x"00000000",
    32433 => x"00000000", 32434 => x"00000000", 32435 => x"00000000",
    32436 => x"00000000", 32437 => x"00000000", 32438 => x"00000000",
    32439 => x"00000000", 32440 => x"00000000", 32441 => x"00000000",
    32442 => x"00000000", 32443 => x"00000000", 32444 => x"00000000",
    32445 => x"00000000", 32446 => x"00000000", 32447 => x"00000000",
    32448 => x"00000000", 32449 => x"00000000", 32450 => x"00000000",
    32451 => x"00000000", 32452 => x"00000000", 32453 => x"00000000",
    32454 => x"00000000", 32455 => x"00000000", 32456 => x"00000000",
    32457 => x"00000000", 32458 => x"00000000", 32459 => x"00000000",
    32460 => x"00000000", 32461 => x"00000000", 32462 => x"00000000",
    32463 => x"00000000", 32464 => x"00000000", 32465 => x"00000000",
    32466 => x"00000000", 32467 => x"00000000", 32468 => x"00000000",
    32469 => x"00000000", 32470 => x"00000000", 32471 => x"00000000",
    32472 => x"00000000", 32473 => x"00000000", 32474 => x"00000000",
    32475 => x"00000000", 32476 => x"00000000", 32477 => x"00000000",
    32478 => x"00000000", 32479 => x"00000000", 32480 => x"00000000",
    32481 => x"00000000", 32482 => x"00000000", 32483 => x"00000000",
    32484 => x"00000000", 32485 => x"00000000", 32486 => x"00000000",
    32487 => x"00000000", 32488 => x"00000000", 32489 => x"00000000",
    32490 => x"00000000", 32491 => x"00000000", 32492 => x"00000000",
    32493 => x"00000000", 32494 => x"00000000", 32495 => x"00000000",
    32496 => x"00000000", 32497 => x"00000000", 32498 => x"00000000",
    32499 => x"00000000", 32500 => x"00000000", 32501 => x"00000000",
    32502 => x"00000000", 32503 => x"00000000", 32504 => x"00000000",
    32505 => x"00000000", 32506 => x"00000000", 32507 => x"00000000",
    32508 => x"00000000", 32509 => x"00000000", 32510 => x"00000000",
    32511 => x"00000000", 32512 => x"00000000", 32513 => x"00000000",
    32514 => x"00000000", 32515 => x"00000000", 32516 => x"00000000",
    32517 => x"00000000", 32518 => x"00000000", 32519 => x"00000000",
    32520 => x"00000000", 32521 => x"00000000", 32522 => x"00000000",
    32523 => x"00000000", 32524 => x"00000000", 32525 => x"00000000",
    32526 => x"00000000", 32527 => x"00000000", 32528 => x"00000000",
    32529 => x"00000000", 32530 => x"00000000", 32531 => x"00000000",
    32532 => x"00000000", 32533 => x"00000000", 32534 => x"00000000",
    32535 => x"00000000", 32536 => x"00000000", 32537 => x"00000000",
    32538 => x"00000000", 32539 => x"00000000", 32540 => x"00000000",
    32541 => x"00000000", 32542 => x"00000000", 32543 => x"00000000",
    32544 => x"00000000", 32545 => x"00000000", 32546 => x"00000000",
    32547 => x"00000000", 32548 => x"00000000", 32549 => x"00000000",
    32550 => x"00000000", 32551 => x"00000000", 32552 => x"00000000",
    32553 => x"00000000", 32554 => x"00000000", 32555 => x"00000000",
    32556 => x"00000000", 32557 => x"00000000", 32558 => x"00000000",
    32559 => x"00000000", 32560 => x"00000000", 32561 => x"00000000",
    32562 => x"00000000", 32563 => x"00000000", 32564 => x"00000000",
    32565 => x"00000000", 32566 => x"00000000", 32567 => x"00000000",
    32568 => x"00000000", 32569 => x"00000000", 32570 => x"00000000",
    32571 => x"00000000", 32572 => x"00000000", 32573 => x"00000000",
    32574 => x"00000000", 32575 => x"00000000", 32576 => x"00000000",
    32577 => x"00000000", 32578 => x"00000000", 32579 => x"00000000",
    32580 => x"00000000", 32581 => x"00000000", 32582 => x"00000000",
    32583 => x"00000000", 32584 => x"00000000", 32585 => x"00000000",
    32586 => x"00000000", 32587 => x"00000000", 32588 => x"00000000",
    32589 => x"00000000", 32590 => x"00000000", 32591 => x"00000000",
    32592 => x"00000000", 32593 => x"00000000", 32594 => x"00000000",
    32595 => x"00000000", 32596 => x"00000000", 32597 => x"00000000",
    32598 => x"00000000", 32599 => x"00000000", 32600 => x"00000000",
    32601 => x"00000000", 32602 => x"00000000", 32603 => x"00000000",
    32604 => x"00000000", 32605 => x"00000000", 32606 => x"00000000",
    32607 => x"00000000", 32608 => x"00000000", 32609 => x"00000000",
    32610 => x"00000000", 32611 => x"00000000", 32612 => x"00000000",
    32613 => x"00000000", 32614 => x"00000000", 32615 => x"00000000",
    32616 => x"00000000", 32617 => x"00000000", 32618 => x"00000000",
    32619 => x"00000000", 32620 => x"00000000", 32621 => x"00000000",
    32622 => x"00000000", 32623 => x"00000000", 32624 => x"00000000",
    32625 => x"00000000", 32626 => x"00000000", 32627 => x"00000000",
    32628 => x"00000000", 32629 => x"00000000", 32630 => x"00000000",
    32631 => x"00000000", 32632 => x"00000000", 32633 => x"00000000",
    32634 => x"00000000", 32635 => x"00000000", 32636 => x"00000000",
    32637 => x"00000000", 32638 => x"00000000", 32639 => x"00000000",
    32640 => x"00000000", 32641 => x"00000000", 32642 => x"00000000",
    32643 => x"00000000", 32644 => x"00000000", 32645 => x"00000000",
    32646 => x"00000000", 32647 => x"00000000", 32648 => x"00000000",
    32649 => x"00000000", 32650 => x"00000000", 32651 => x"00000000",
    32652 => x"00000000", 32653 => x"00000000", 32654 => x"00000000",
    32655 => x"00000000", 32656 => x"00000000", 32657 => x"00000000",
    32658 => x"00000000", 32659 => x"00000000", 32660 => x"00000000",
    32661 => x"00000000", 32662 => x"00000000", 32663 => x"00000000",
    32664 => x"00000000", 32665 => x"00000000", 32666 => x"00000000",
    32667 => x"00000000", 32668 => x"00000000", 32669 => x"00000000",
    32670 => x"00000000", 32671 => x"00000000", 32672 => x"00000000",
    32673 => x"00000000", 32674 => x"00000000", 32675 => x"00000000",
    32676 => x"00000000", 32677 => x"00000000", 32678 => x"00000000",
    32679 => x"00000000", 32680 => x"00000000", 32681 => x"00000000",
    32682 => x"00000000", 32683 => x"00000000", 32684 => x"00000000",
    32685 => x"00000000", 32686 => x"00000000", 32687 => x"00000000",
    32688 => x"00000000", 32689 => x"00000000", 32690 => x"00000000",
    32691 => x"00000000", 32692 => x"00000000", 32693 => x"00000000",
    32694 => x"00000000", 32695 => x"00000000", 32696 => x"00000000",
    32697 => x"00000000", 32698 => x"00000000", 32699 => x"00000000",
    32700 => x"00000000", 32701 => x"00000000", 32702 => x"00000000",
    32703 => x"00000000", 32704 => x"00000000", 32705 => x"00000000",
    32706 => x"00000000", 32707 => x"00000000", 32708 => x"00000000",
    32709 => x"00000000", 32710 => x"00000000", 32711 => x"00000000",
    32712 => x"00000000", 32713 => x"00000000", 32714 => x"00000000",
    32715 => x"00000000", 32716 => x"00000000", 32717 => x"00000000",
    32718 => x"00000000", 32719 => x"00000000", 32720 => x"00000000",
    32721 => x"00000000", 32722 => x"00000000", 32723 => x"00000000",
    32724 => x"00000000", 32725 => x"00000000", 32726 => x"00000000",
    32727 => x"00000000", 32728 => x"00000000", 32729 => x"00000000",
    32730 => x"00000000", 32731 => x"00000000", 32732 => x"00000000",
    32733 => x"00000000", 32734 => x"00000000", 32735 => x"00000000",
    32736 => x"00000000", 32737 => x"00000000", 32738 => x"00000000",
    32739 => x"00000000", 32740 => x"00000000", 32741 => x"00000000",
    32742 => x"00000000", 32743 => x"00000000", 32744 => x"00000000",
    32745 => x"00000000", 32746 => x"00000000", 32747 => x"00000000",
    32748 => x"00000000", 32749 => x"00000000", 32750 => x"00000000",
    32751 => x"00000000", 32752 => x"00000000", 32753 => x"00000000",
    32754 => x"00000000", 32755 => x"00000000", 32756 => x"00000000",
    32757 => x"00000000", 32758 => x"00000000", 32759 => x"00000000",
    32760 => x"00000000", 32761 => x"00000000", 32762 => x"00000000",
    32763 => x"00000000", 32764 => x"00000000", 32765 => x"00000000",
    32766 => x"00000000", 32767 => x"00000000");
end wrc_bin_pkg;
